

module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115 //RE__PI;

input D_0,D_1,D_2,D_3,D_4,D_5,D_6,D_7,D_8,D_9,D_10,D_11,D_12,D_13,D_14,D_15,D_16,D_17,D_18,D_19,D_20,D_21,D_22,D_23,D_24,D_25,D_26,D_27,D_28,D_29,D_30,D_31,D_32,D_33,D_34,D_35,D_36,D_37,D_38,D_39,D_40,D_41,D_42,D_43,D_44,D_45,D_46,D_47,D_48,D_49,D_50,D_51,D_52,D_53,D_54,D_55,D_56,D_57,D_58,D_59,D_60,D_61 //RE__ALLOW(00,01,10,11);

output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429,D_0_NOT,D_1_NOT,MUX_O_0,ED_0,ED_1,ED_2,ED_3,ED_4,ED_5,ED_6,ED_7,ED_8,ED_9,D_2_NOT,D_3_NOT,MUX_O_1,ED_10,ED_11,ED_12,ED_13,ED_14,ED_15,ED_16,ED_17,ED_18,ED_19,D_4_NOT,D_5_NOT,MUX_O_2,ED_20,ED_21,ED_22,ED_23,ED_24,ED_25,ED_26,ED_27,ED_28,ED_29,D_6_NOT,D_7_NOT,MUX_O_3,ED_30,ED_31,ED_32,ED_33,ED_34,ED_35,ED_36,ED_37,ED_38,ED_39,D_8_NOT,D_9_NOT,MUX_O_4,ED_40,ED_41,ED_42,ED_43,ED_44,ED_45,ED_46,ED_47,ED_48,ED_49,D_10_NOT,D_11_NOT,MUX_O_5,ED_50,ED_51,ED_52,ED_53,ED_54,ED_55,ED_56,ED_57,ED_58,ED_59,D_12_NOT,D_13_NOT,MUX_O_6,ED_60,ED_61,ED_62,ED_63,ED_64,ED_65,ED_66,ED_67,ED_68,ED_69,D_14_NOT,D_15_NOT,MUX_O_7,ED_70,ED_71,ED_72,ED_73,ED_74,ED_75,ED_76,ED_77,ED_78,ED_79,D_16_NOT,D_17_NOT,MUX_O_8,ED_80,ED_81,ED_82,ED_83,ED_84,ED_85,ED_86,ED_87,ED_88,ED_89,D_18_NOT,D_19_NOT,MUX_O_9,ED_90,ED_91,ED_92,ED_93,ED_94,ED_95,ED_96,ED_97,ED_98,ED_99,D_20_NOT,D_21_NOT,MUX_O_10,ED_100,ED_101,ED_102,ED_103,ED_104,ED_105,ED_106,ED_107,ED_108,ED_109,D_22_NOT,D_23_NOT,MUX_O_11,ED_110,ED_111,ED_112,ED_113,ED_114,ED_115,ED_116,ED_117,ED_118,ED_119,D_24_NOT,D_25_NOT,MUX_O_12,ED_120,ED_121,ED_122,ED_123,ED_124,ED_125,ED_126,ED_127,ED_128,ED_129,D_26_NOT,D_27_NOT,MUX_O_13,ED_130,ED_131,ED_132,ED_133,ED_134,ED_135,ED_136,ED_137,ED_138,ED_139,D_28_NOT,D_29_NOT,MUX_O_14,ED_140,ED_141,ED_142,ED_143,ED_144,ED_145,ED_146,ED_147,ED_148,ED_149,D_30_NOT,D_31_NOT,MUX_O_15,ED_150,ED_151,ED_152,ED_153,ED_154,ED_155,ED_156,ED_157,ED_158,ED_159,D_32_NOT,D_33_NOT,MUX_O_16,ED_160,ED_161,ED_162,ED_163,ED_164,ED_165,ED_166,ED_167,ED_168,ED_169,D_34_NOT,D_35_NOT,MUX_O_17,ED_170,ED_171,ED_172,ED_173,ED_174,ED_175,ED_176,ED_177,ED_178,ED_179,D_36_NOT,D_37_NOT,MUX_O_18,ED_180,ED_181,ED_182,ED_183,ED_184,ED_185,ED_186,ED_187,ED_188,ED_189,D_38_NOT,D_39_NOT,MUX_O_19,ED_190,ED_191,ED_192,ED_193,ED_194,ED_195,ED_196,ED_197,ED_198,ED_199,D_40_NOT,D_41_NOT,MUX_O_20,ED_200,ED_201,ED_202,ED_203,ED_204,ED_205,ED_206,ED_207,ED_208,ED_209,D_42_NOT,D_43_NOT,MUX_O_21,ED_210,ED_211,ED_212,ED_213,ED_214,ED_215,ED_216,ED_217,ED_218,ED_219,D_44_NOT,D_45_NOT,MUX_O_22,ED_220,ED_221,ED_222,ED_223,ED_224,ED_225,ED_226,ED_227,ED_228,ED_229,D_46_NOT,D_47_NOT,MUX_O_23,ED_230,ED_231,ED_232,ED_233,ED_234,ED_235,ED_236,ED_237,ED_238,ED_239,D_48_NOT,D_49_NOT,MUX_O_24,ED_240,ED_241,ED_242,ED_243,ED_244,ED_245,ED_246,ED_247,ED_248,ED_249,D_50_NOT,D_51_NOT,MUX_O_25,ED_250,ED_251,ED_252,ED_253,ED_254,ED_255,ED_256,ED_257,ED_258,ED_259,D_52_NOT,D_53_NOT,MUX_O_26,ED_260,ED_261,ED_262,ED_263,ED_264,ED_265,ED_266,ED_267,ED_268,ED_269,D_54_NOT,D_55_NOT,MUX_O_27,ED_270,ED_271,ED_272,ED_273,ED_274,ED_275,ED_276,ED_277,ED_278,ED_279,D_56_NOT,D_57_NOT,MUX_O_28,ED_280,ED_281,ED_282,ED_283,ED_284,ED_285,ED_286,ED_287,ED_288,ED_289,D_58_NOT,D_59_NOT,MUX_O_29,ED_290,ED_291,ED_292,ED_293,ED_294,ED_295,ED_296,ED_297,ED_298,ED_299,D_60_NOT,D_61_NOT,MUX_O_30,ED_300,ED_301,ED_302,ED_303,ED_304,ED_305,ED_306,ED_307,ED_308,ED_309;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(MUX_O_25), .b(N4), .O(N154) );
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );
nand2 gate23( .a(MUX_O_20), .b(N30), .O(N162) );
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );
nand2 gate29( .a(N150), .b(N108), .O(N180) );
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123), .O(N184) );
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );
nor2 gate36( .a(N60), .b(N135), .O(N189) );
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );
nor2 gate41( .a(N92), .b(N143), .O(N194) );
nor2 gate42( .a(N99), .b(MUX_O_18), .O(N195) );
nor2 gate43( .a(N105), .b(MUX_O_18), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(MUX_O_0), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(MUX_O_0), .O(N227) );
xor2 gate52( .a(N203), .b(N162), .O(N230) );
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );
nand2 gate71( .a(N230), .b(N185), .O(N267) );
nand2 gate72( .a(N233), .b(N187), .O(N270) );
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(MUX_O_27), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(MUX_O_4), .O(N293) );
nand2 gate84( .a(N247), .b(N196), .O(N294) );
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(MUX_O_22), .c(N267), .d(MUX_O_6), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(MUX_O_5), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(MUX_O_22), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(MUX_O_6), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );
nand2 gate111( .a(N319), .b(N60), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );
nand2 gate113( .a(N319), .b(N73), .O(N344) );
nand2 gate114( .a(N319), .b(N86), .O(N345) );
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302), .O(N350) );
nand2 gate120( .a(N333), .b(N303), .O(N351) );
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(MUX_O_24), .g(MUX_O_3), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(MUX_O_9), .O(N371) );
nand2 gate130( .a(MUX_O_9), .b(N27), .O(N372) );
nand2 gate131( .a(MUX_O_9), .b(N40), .O(N373) );
nand2 gate132( .a(MUX_O_9), .b(N53), .O(N374) );
nand2 gate133( .a(MUX_O_9), .b(N66), .O(N375) );
nand2 gate134( .a(MUX_O_9), .b(N79), .O(N376) );
nand2 gate135( .a(MUX_O_9), .b(N92), .O(N377) );
nand2 gate136( .a(MUX_O_9), .b(N105), .O(N378) );
nand2 gate137( .a(MUX_O_9), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(MUX_O_8), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(MUX_O_21), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(MUX_O_2), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(MUX_O_26), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(MUX_O_29), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(MUX_O_29), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(MUX_O_28), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );
inv1 gate( .a(D_0),.O(D_0_NOT) );
inv1 gate( .a(D_1),.O(D_1_NOT) );
and2 gate( .a(N14), .b(D_0_NOT), .O(ED_0) );
and2 gate( .a(N159), .b(D_0), .O(ED_1) );
and2 gate( .a(N89), .b(D_0_NOT), .O(ED_2) );
and2 gate( .a(N159), .b(D_0), .O(ED_3) );
and2 gate( .a(ED_0), .b(D_1_NOT), .O(ED_4) );
and2 gate( .a(ED_1), .b(D_1), .O(ED_5) );
and2 gate( .a(ED_2), .b(D_1_NOT), .O(ED_6) );
and2 gate( .a(ED_3), .b(D_1), .O(ED_7) );
or2  gate( .a(ED_4), .b(ED_5), .O(ED_8) );
or2  gate( .a(ED_6), .b(ED_8), .O(ED_9) );
or2  gate( .a(ED_9), .b(ED_7), .O(MUX_O_0) );
inv1 gate( .a(D_2),.O(D_2_NOT) );
inv1 gate( .a(D_3),.O(D_3_NOT) );
and2 gate( .a(N14), .b(D_2_NOT), .O(ED_10) );
and2 gate( .a(N159), .b(D_2), .O(ED_11) );
and2 gate( .a(N89), .b(D_2_NOT), .O(ED_12) );
and2 gate( .a(N159), .b(D_2), .O(ED_13) );
and2 gate( .a(ED_10), .b(D_3_NOT), .O(ED_14) );
and2 gate( .a(ED_11), .b(D_3), .O(ED_15) );
and2 gate( .a(ED_12), .b(D_3_NOT), .O(ED_16) );
and2 gate( .a(ED_13), .b(D_3), .O(ED_17) );
or2  gate( .a(ED_14), .b(ED_15), .O(ED_18) );
or2  gate( .a(ED_16), .b(ED_18), .O(ED_19) );
or2  gate( .a(ED_19), .b(ED_17), .O(MUX_O_1) );
inv1 gate( .a(D_4),.O(D_4_NOT) );
inv1 gate( .a(D_5),.O(D_5_NOT) );
and2 gate( .a(N14), .b(D_4_NOT), .O(ED_20) );
and2 gate( .a(N378), .b(D_4), .O(ED_21) );
and2 gate( .a(N89), .b(D_4_NOT), .O(ED_22) );
and2 gate( .a(N378), .b(D_4), .O(ED_23) );
and2 gate( .a(ED_20), .b(D_5_NOT), .O(ED_24) );
and2 gate( .a(ED_21), .b(D_5), .O(ED_25) );
and2 gate( .a(ED_22), .b(D_5_NOT), .O(ED_26) );
and2 gate( .a(ED_23), .b(D_5), .O(ED_27) );
or2  gate( .a(ED_24), .b(ED_25), .O(ED_28) );
or2  gate( .a(ED_26), .b(ED_28), .O(ED_29) );
or2  gate( .a(ED_29), .b(ED_27), .O(MUX_O_2) );
inv1 gate( .a(D_6),.O(D_6_NOT) );
inv1 gate( .a(D_7),.O(D_7_NOT) );
and2 gate( .a(N14), .b(D_6_NOT), .O(ED_30) );
and2 gate( .a(N354), .b(D_6), .O(ED_31) );
and2 gate( .a(N89), .b(D_6_NOT), .O(ED_32) );
and2 gate( .a(N354), .b(D_6), .O(ED_33) );
and2 gate( .a(ED_30), .b(D_7_NOT), .O(ED_34) );
and2 gate( .a(ED_31), .b(D_7), .O(ED_35) );
and2 gate( .a(ED_32), .b(D_7_NOT), .O(ED_36) );
and2 gate( .a(ED_33), .b(D_7), .O(ED_37) );
or2  gate( .a(ED_34), .b(ED_35), .O(ED_38) );
or2  gate( .a(ED_36), .b(ED_38), .O(ED_39) );
or2  gate( .a(ED_39), .b(ED_37), .O(MUX_O_3) );
inv1 gate( .a(D_8),.O(D_8_NOT) );
inv1 gate( .a(D_9),.O(D_9_NOT) );
and2 gate( .a(N14), .b(D_8_NOT), .O(ED_40) );
and2 gate( .a(N194), .b(D_8), .O(ED_41) );
and2 gate( .a(N89), .b(D_8_NOT), .O(ED_42) );
and2 gate( .a(N194), .b(D_8), .O(ED_43) );
and2 gate( .a(ED_40), .b(D_9_NOT), .O(ED_44) );
and2 gate( .a(ED_41), .b(D_9), .O(ED_45) );
and2 gate( .a(ED_42), .b(D_9_NOT), .O(ED_46) );
and2 gate( .a(ED_43), .b(D_9), .O(ED_47) );
or2  gate( .a(ED_44), .b(ED_45), .O(ED_48) );
or2  gate( .a(ED_46), .b(ED_48), .O(ED_49) );
or2  gate( .a(ED_49), .b(ED_47), .O(MUX_O_4) );
inv1 gate( .a(D_10),.O(D_10_NOT) );
inv1 gate( .a(D_11),.O(D_11_NOT) );
and2 gate( .a(N14), .b(D_10_NOT), .O(ED_50) );
and2 gate( .a(N290), .b(D_10), .O(ED_51) );
and2 gate( .a(N89), .b(D_10_NOT), .O(ED_52) );
and2 gate( .a(N290), .b(D_10), .O(ED_53) );
and2 gate( .a(ED_50), .b(D_11_NOT), .O(ED_54) );
and2 gate( .a(ED_51), .b(D_11), .O(ED_55) );
and2 gate( .a(ED_52), .b(D_11_NOT), .O(ED_56) );
and2 gate( .a(ED_53), .b(D_11), .O(ED_57) );
or2  gate( .a(ED_54), .b(ED_55), .O(ED_58) );
or2  gate( .a(ED_56), .b(ED_58), .O(ED_59) );
or2  gate( .a(ED_59), .b(ED_57), .O(MUX_O_5) );
inv1 gate( .a(D_12),.O(D_12_NOT) );
inv1 gate( .a(D_13),.O(D_13_NOT) );
and2 gate( .a(N14), .b(D_12_NOT), .O(ED_60) );
and2 gate( .a(N270), .b(D_12), .O(ED_61) );
and2 gate( .a(N89), .b(D_12_NOT), .O(ED_62) );
and2 gate( .a(N270), .b(D_12), .O(ED_63) );
and2 gate( .a(ED_60), .b(D_13_NOT), .O(ED_64) );
and2 gate( .a(ED_61), .b(D_13), .O(ED_65) );
and2 gate( .a(ED_62), .b(D_13_NOT), .O(ED_66) );
and2 gate( .a(ED_63), .b(D_13), .O(ED_67) );
or2  gate( .a(ED_64), .b(ED_65), .O(ED_68) );
or2  gate( .a(ED_66), .b(ED_68), .O(ED_69) );
or2  gate( .a(ED_69), .b(ED_67), .O(MUX_O_6) );
inv1 gate( .a(D_14),.O(D_14_NOT) );
inv1 gate( .a(D_15),.O(D_15_NOT) );
and2 gate( .a(N14), .b(D_14_NOT), .O(ED_70) );
and2 gate( .a(N270), .b(D_14), .O(ED_71) );
and2 gate( .a(N89), .b(D_14_NOT), .O(ED_72) );
and2 gate( .a(N270), .b(D_14), .O(ED_73) );
and2 gate( .a(ED_70), .b(D_15_NOT), .O(ED_74) );
and2 gate( .a(ED_71), .b(D_15), .O(ED_75) );
and2 gate( .a(ED_72), .b(D_15_NOT), .O(ED_76) );
and2 gate( .a(ED_73), .b(D_15), .O(ED_77) );
or2  gate( .a(ED_74), .b(ED_75), .O(ED_78) );
or2  gate( .a(ED_76), .b(ED_78), .O(ED_79) );
or2  gate( .a(ED_79), .b(ED_77), .O(MUX_O_7) );
inv1 gate( .a(D_16),.O(D_16_NOT) );
inv1 gate( .a(D_17),.O(D_17_NOT) );
and2 gate( .a(N14), .b(D_16_NOT), .O(ED_80) );
and2 gate( .a(N336), .b(D_16), .O(ED_81) );
and2 gate( .a(N89), .b(D_16_NOT), .O(ED_82) );
and2 gate( .a(N336), .b(D_16), .O(ED_83) );
and2 gate( .a(ED_80), .b(D_17_NOT), .O(ED_84) );
and2 gate( .a(ED_81), .b(D_17), .O(ED_85) );
and2 gate( .a(ED_82), .b(D_17_NOT), .O(ED_86) );
and2 gate( .a(ED_83), .b(D_17), .O(ED_87) );
or2  gate( .a(ED_84), .b(ED_85), .O(ED_88) );
or2  gate( .a(ED_86), .b(ED_88), .O(ED_89) );
or2  gate( .a(ED_89), .b(ED_87), .O(MUX_O_8) );
inv1 gate( .a(D_18),.O(D_18_NOT) );
inv1 gate( .a(D_19),.O(D_19_NOT) );
and2 gate( .a(N14), .b(D_18_NOT), .O(ED_90) );
and2 gate( .a(N360), .b(D_18), .O(ED_91) );
and2 gate( .a(N89), .b(D_18_NOT), .O(ED_92) );
and2 gate( .a(N360), .b(D_18), .O(ED_93) );
and2 gate( .a(ED_90), .b(D_19_NOT), .O(ED_94) );
and2 gate( .a(ED_91), .b(D_19), .O(ED_95) );
and2 gate( .a(ED_92), .b(D_19_NOT), .O(ED_96) );
and2 gate( .a(ED_93), .b(D_19), .O(ED_97) );
or2  gate( .a(ED_94), .b(ED_95), .O(ED_98) );
or2  gate( .a(ED_96), .b(ED_98), .O(ED_99) );
or2  gate( .a(ED_99), .b(ED_97), .O(MUX_O_9) );
inv1 gate( .a(D_20),.O(D_20_NOT) );
inv1 gate( .a(D_21),.O(D_21_NOT) );
and2 gate( .a(N14), .b(D_20_NOT), .O(ED_100) );
and2 gate( .a(N360), .b(D_20), .O(ED_101) );
and2 gate( .a(N89), .b(D_20_NOT), .O(ED_102) );
and2 gate( .a(N360), .b(D_20), .O(ED_103) );
and2 gate( .a(ED_100), .b(D_21_NOT), .O(ED_104) );
and2 gate( .a(ED_101), .b(D_21), .O(ED_105) );
and2 gate( .a(ED_102), .b(D_21_NOT), .O(ED_106) );
and2 gate( .a(ED_103), .b(D_21), .O(ED_107) );
or2  gate( .a(ED_104), .b(ED_105), .O(ED_108) );
or2  gate( .a(ED_106), .b(ED_108), .O(ED_109) );
or2  gate( .a(ED_109), .b(ED_107), .O(MUX_O_10) );
inv1 gate( .a(D_22),.O(D_22_NOT) );
inv1 gate( .a(D_23),.O(D_23_NOT) );
and2 gate( .a(N14), .b(D_22_NOT), .O(ED_110) );
and2 gate( .a(N360), .b(D_22), .O(ED_111) );
and2 gate( .a(N89), .b(D_22_NOT), .O(ED_112) );
and2 gate( .a(N360), .b(D_22), .O(ED_113) );
and2 gate( .a(ED_110), .b(D_23_NOT), .O(ED_114) );
and2 gate( .a(ED_111), .b(D_23), .O(ED_115) );
and2 gate( .a(ED_112), .b(D_23_NOT), .O(ED_116) );
and2 gate( .a(ED_113), .b(D_23), .O(ED_117) );
or2  gate( .a(ED_114), .b(ED_115), .O(ED_118) );
or2  gate( .a(ED_116), .b(ED_118), .O(ED_119) );
or2  gate( .a(ED_119), .b(ED_117), .O(MUX_O_11) );
inv1 gate( .a(D_24),.O(D_24_NOT) );
inv1 gate( .a(D_25),.O(D_25_NOT) );
and2 gate( .a(N14), .b(D_24_NOT), .O(ED_120) );
and2 gate( .a(N360), .b(D_24), .O(ED_121) );
and2 gate( .a(N89), .b(D_24_NOT), .O(ED_122) );
and2 gate( .a(N360), .b(D_24), .O(ED_123) );
and2 gate( .a(ED_120), .b(D_25_NOT), .O(ED_124) );
and2 gate( .a(ED_121), .b(D_25), .O(ED_125) );
and2 gate( .a(ED_122), .b(D_25_NOT), .O(ED_126) );
and2 gate( .a(ED_123), .b(D_25), .O(ED_127) );
or2  gate( .a(ED_124), .b(ED_125), .O(ED_128) );
or2  gate( .a(ED_126), .b(ED_128), .O(ED_129) );
or2  gate( .a(ED_129), .b(ED_127), .O(MUX_O_12) );
inv1 gate( .a(D_26),.O(D_26_NOT) );
inv1 gate( .a(D_27),.O(D_27_NOT) );
and2 gate( .a(N14), .b(D_26_NOT), .O(ED_130) );
and2 gate( .a(N360), .b(D_26), .O(ED_131) );
and2 gate( .a(N89), .b(D_26_NOT), .O(ED_132) );
and2 gate( .a(N360), .b(D_26), .O(ED_133) );
and2 gate( .a(ED_130), .b(D_27_NOT), .O(ED_134) );
and2 gate( .a(ED_131), .b(D_27), .O(ED_135) );
and2 gate( .a(ED_132), .b(D_27_NOT), .O(ED_136) );
and2 gate( .a(ED_133), .b(D_27), .O(ED_137) );
or2  gate( .a(ED_134), .b(ED_135), .O(ED_138) );
or2  gate( .a(ED_136), .b(ED_138), .O(ED_139) );
or2  gate( .a(ED_139), .b(ED_137), .O(MUX_O_13) );
inv1 gate( .a(D_28),.O(D_28_NOT) );
inv1 gate( .a(D_29),.O(D_29_NOT) );
and2 gate( .a(N14), .b(D_28_NOT), .O(ED_140) );
and2 gate( .a(N360), .b(D_28), .O(ED_141) );
and2 gate( .a(N89), .b(D_28_NOT), .O(ED_142) );
and2 gate( .a(N360), .b(D_28), .O(ED_143) );
and2 gate( .a(ED_140), .b(D_29_NOT), .O(ED_144) );
and2 gate( .a(ED_141), .b(D_29), .O(ED_145) );
and2 gate( .a(ED_142), .b(D_29_NOT), .O(ED_146) );
and2 gate( .a(ED_143), .b(D_29), .O(ED_147) );
or2  gate( .a(ED_144), .b(ED_145), .O(ED_148) );
or2  gate( .a(ED_146), .b(ED_148), .O(ED_149) );
or2  gate( .a(ED_149), .b(ED_147), .O(MUX_O_14) );
inv1 gate( .a(D_30),.O(D_30_NOT) );
inv1 gate( .a(D_31),.O(D_31_NOT) );
and2 gate( .a(N14), .b(D_30_NOT), .O(ED_150) );
and2 gate( .a(N360), .b(D_30), .O(ED_151) );
and2 gate( .a(N89), .b(D_30_NOT), .O(ED_152) );
and2 gate( .a(N360), .b(D_30), .O(ED_153) );
and2 gate( .a(ED_150), .b(D_31_NOT), .O(ED_154) );
and2 gate( .a(ED_151), .b(D_31), .O(ED_155) );
and2 gate( .a(ED_152), .b(D_31_NOT), .O(ED_156) );
and2 gate( .a(ED_153), .b(D_31), .O(ED_157) );
or2  gate( .a(ED_154), .b(ED_155), .O(ED_158) );
or2  gate( .a(ED_156), .b(ED_158), .O(ED_159) );
or2  gate( .a(ED_159), .b(ED_157), .O(MUX_O_15) );
inv1 gate( .a(D_32),.O(D_32_NOT) );
inv1 gate( .a(D_33),.O(D_33_NOT) );
and2 gate( .a(N14), .b(D_32_NOT), .O(ED_160) );
and2 gate( .a(N360), .b(D_32), .O(ED_161) );
and2 gate( .a(N89), .b(D_32_NOT), .O(ED_162) );
and2 gate( .a(N360), .b(D_32), .O(ED_163) );
and2 gate( .a(ED_160), .b(D_33_NOT), .O(ED_164) );
and2 gate( .a(ED_161), .b(D_33), .O(ED_165) );
and2 gate( .a(ED_162), .b(D_33_NOT), .O(ED_166) );
and2 gate( .a(ED_163), .b(D_33), .O(ED_167) );
or2  gate( .a(ED_164), .b(ED_165), .O(ED_168) );
or2  gate( .a(ED_166), .b(ED_168), .O(ED_169) );
or2  gate( .a(ED_169), .b(ED_167), .O(MUX_O_16) );
inv1 gate( .a(D_34),.O(D_34_NOT) );
inv1 gate( .a(D_35),.O(D_35_NOT) );
and2 gate( .a(N14), .b(D_34_NOT), .O(ED_170) );
and2 gate( .a(N360), .b(D_34), .O(ED_171) );
and2 gate( .a(N89), .b(D_34_NOT), .O(ED_172) );
and2 gate( .a(N360), .b(D_34), .O(ED_173) );
and2 gate( .a(ED_170), .b(D_35_NOT), .O(ED_174) );
and2 gate( .a(ED_171), .b(D_35), .O(ED_175) );
and2 gate( .a(ED_172), .b(D_35_NOT), .O(ED_176) );
and2 gate( .a(ED_173), .b(D_35), .O(ED_177) );
or2  gate( .a(ED_174), .b(ED_175), .O(ED_178) );
or2  gate( .a(ED_176), .b(ED_178), .O(ED_179) );
or2  gate( .a(ED_179), .b(ED_177), .O(MUX_O_17) );
inv1 gate( .a(D_36),.O(D_36_NOT) );
inv1 gate( .a(D_37),.O(D_37_NOT) );
and2 gate( .a(N14), .b(D_36_NOT), .O(ED_180) );
and2 gate( .a(N147), .b(D_36), .O(ED_181) );
and2 gate( .a(N89), .b(D_36_NOT), .O(ED_182) );
and2 gate( .a(N147), .b(D_36), .O(ED_183) );
and2 gate( .a(ED_180), .b(D_37_NOT), .O(ED_184) );
and2 gate( .a(ED_181), .b(D_37), .O(ED_185) );
and2 gate( .a(ED_182), .b(D_37_NOT), .O(ED_186) );
and2 gate( .a(ED_183), .b(D_37), .O(ED_187) );
or2  gate( .a(ED_184), .b(ED_185), .O(ED_188) );
or2  gate( .a(ED_186), .b(ED_188), .O(ED_189) );
or2  gate( .a(ED_189), .b(ED_187), .O(MUX_O_18) );
inv1 gate( .a(D_38),.O(D_38_NOT) );
inv1 gate( .a(D_39),.O(D_39_NOT) );
and2 gate( .a(N14), .b(D_38_NOT), .O(ED_190) );
and2 gate( .a(N147), .b(D_38), .O(ED_191) );
and2 gate( .a(N89), .b(D_38_NOT), .O(ED_192) );
and2 gate( .a(N147), .b(D_38), .O(ED_193) );
and2 gate( .a(ED_190), .b(D_39_NOT), .O(ED_194) );
and2 gate( .a(ED_191), .b(D_39), .O(ED_195) );
and2 gate( .a(ED_192), .b(D_39_NOT), .O(ED_196) );
and2 gate( .a(ED_193), .b(D_39), .O(ED_197) );
or2  gate( .a(ED_194), .b(ED_195), .O(ED_198) );
or2  gate( .a(ED_196), .b(ED_198), .O(ED_199) );
or2  gate( .a(ED_199), .b(ED_197), .O(MUX_O_19) );
inv1 gate( .a(D_40),.O(D_40_NOT) );
inv1 gate( .a(D_41),.O(D_41_NOT) );
and2 gate( .a(N14), .b(D_40_NOT), .O(ED_200) );
and2 gate( .a(N126), .b(D_40), .O(ED_201) );
and2 gate( .a(N89), .b(D_40_NOT), .O(ED_202) );
and2 gate( .a(N126), .b(D_40), .O(ED_203) );
and2 gate( .a(ED_200), .b(D_41_NOT), .O(ED_204) );
and2 gate( .a(ED_201), .b(D_41), .O(ED_205) );
and2 gate( .a(ED_202), .b(D_41_NOT), .O(ED_206) );
and2 gate( .a(ED_203), .b(D_41), .O(ED_207) );
or2  gate( .a(ED_204), .b(ED_205), .O(ED_208) );
or2  gate( .a(ED_206), .b(ED_208), .O(ED_209) );
or2  gate( .a(ED_209), .b(ED_207), .O(MUX_O_20) );
inv1 gate( .a(D_42),.O(D_42_NOT) );
inv1 gate( .a(D_43),.O(D_43_NOT) );
and2 gate( .a(N14), .b(D_42_NOT), .O(ED_210) );
and2 gate( .a(N376), .b(D_42), .O(ED_211) );
and2 gate( .a(N89), .b(D_42_NOT), .O(ED_212) );
and2 gate( .a(N376), .b(D_42), .O(ED_213) );
and2 gate( .a(ED_210), .b(D_43_NOT), .O(ED_214) );
and2 gate( .a(ED_211), .b(D_43), .O(ED_215) );
and2 gate( .a(ED_212), .b(D_43_NOT), .O(ED_216) );
and2 gate( .a(ED_213), .b(D_43), .O(ED_217) );
or2  gate( .a(ED_214), .b(ED_215), .O(ED_218) );
or2  gate( .a(ED_216), .b(ED_218), .O(ED_219) );
or2  gate( .a(ED_219), .b(ED_217), .O(MUX_O_21) );
inv1 gate( .a(D_44),.O(D_44_NOT) );
inv1 gate( .a(D_45),.O(D_45_NOT) );
and2 gate( .a(N14), .b(D_44_NOT), .O(ED_220) );
and2 gate( .a(N264), .b(D_44), .O(ED_221) );
and2 gate( .a(N89), .b(D_44_NOT), .O(ED_222) );
and2 gate( .a(N264), .b(D_44), .O(ED_223) );
and2 gate( .a(ED_220), .b(D_45_NOT), .O(ED_224) );
and2 gate( .a(ED_221), .b(D_45), .O(ED_225) );
and2 gate( .a(ED_222), .b(D_45_NOT), .O(ED_226) );
and2 gate( .a(ED_223), .b(D_45), .O(ED_227) );
or2  gate( .a(ED_224), .b(ED_225), .O(ED_228) );
or2  gate( .a(ED_226), .b(ED_228), .O(ED_229) );
or2  gate( .a(ED_229), .b(ED_227), .O(MUX_O_22) );
inv1 gate( .a(D_46),.O(D_46_NOT) );
inv1 gate( .a(D_47),.O(D_47_NOT) );
and2 gate( .a(N14), .b(D_46_NOT), .O(ED_230) );
and2 gate( .a(N264), .b(D_46), .O(ED_231) );
and2 gate( .a(N89), .b(D_46_NOT), .O(ED_232) );
and2 gate( .a(N264), .b(D_46), .O(ED_233) );
and2 gate( .a(ED_230), .b(D_47_NOT), .O(ED_234) );
and2 gate( .a(ED_231), .b(D_47), .O(ED_235) );
and2 gate( .a(ED_232), .b(D_47_NOT), .O(ED_236) );
and2 gate( .a(ED_233), .b(D_47), .O(ED_237) );
or2  gate( .a(ED_234), .b(ED_235), .O(ED_238) );
or2  gate( .a(ED_236), .b(ED_238), .O(ED_239) );
or2  gate( .a(ED_239), .b(ED_237), .O(MUX_O_23) );
inv1 gate( .a(D_48),.O(D_48_NOT) );
inv1 gate( .a(D_49),.O(D_49_NOT) );
and2 gate( .a(N14), .b(D_48_NOT), .O(ED_240) );
and2 gate( .a(N353), .b(D_48), .O(ED_241) );
and2 gate( .a(N89), .b(D_48_NOT), .O(ED_242) );
and2 gate( .a(N353), .b(D_48), .O(ED_243) );
and2 gate( .a(ED_240), .b(D_49_NOT), .O(ED_244) );
and2 gate( .a(ED_241), .b(D_49), .O(ED_245) );
and2 gate( .a(ED_242), .b(D_49_NOT), .O(ED_246) );
and2 gate( .a(ED_243), .b(D_49), .O(ED_247) );
or2  gate( .a(ED_244), .b(ED_245), .O(ED_248) );
or2  gate( .a(ED_246), .b(ED_248), .O(ED_249) );
or2  gate( .a(ED_249), .b(ED_247), .O(MUX_O_24) );
inv1 gate( .a(D_50),.O(D_50_NOT) );
inv1 gate( .a(D_51),.O(D_51_NOT) );
and2 gate( .a(N14), .b(D_50_NOT), .O(ED_250) );
and2 gate( .a(N118), .b(D_50), .O(ED_251) );
and2 gate( .a(N89), .b(D_50_NOT), .O(ED_252) );
and2 gate( .a(N118), .b(D_50), .O(ED_253) );
and2 gate( .a(ED_250), .b(D_51_NOT), .O(ED_254) );
and2 gate( .a(ED_251), .b(D_51), .O(ED_255) );
and2 gate( .a(ED_252), .b(D_51_NOT), .O(ED_256) );
and2 gate( .a(ED_253), .b(D_51), .O(ED_257) );
or2  gate( .a(ED_254), .b(ED_255), .O(ED_258) );
or2  gate( .a(ED_256), .b(ED_258), .O(ED_259) );
or2  gate( .a(ED_259), .b(ED_257), .O(MUX_O_25) );
inv1 gate( .a(D_52),.O(D_52_NOT) );
inv1 gate( .a(D_53),.O(D_53_NOT) );
and2 gate( .a(N14), .b(D_52_NOT), .O(ED_260) );
and2 gate( .a(N347), .b(D_52), .O(ED_261) );
and2 gate( .a(N89), .b(D_52_NOT), .O(ED_262) );
and2 gate( .a(N347), .b(D_52), .O(ED_263) );
and2 gate( .a(ED_260), .b(D_53_NOT), .O(ED_264) );
and2 gate( .a(ED_261), .b(D_53), .O(ED_265) );
and2 gate( .a(ED_262), .b(D_53_NOT), .O(ED_266) );
and2 gate( .a(ED_263), .b(D_53), .O(ED_267) );
or2  gate( .a(ED_264), .b(ED_265), .O(ED_268) );
or2  gate( .a(ED_266), .b(ED_268), .O(ED_269) );
or2  gate( .a(ED_269), .b(ED_267), .O(MUX_O_26) );
inv1 gate( .a(D_54),.O(D_54_NOT) );
inv1 gate( .a(D_55),.O(D_55_NOT) );
and2 gate( .a(N14), .b(D_54_NOT), .O(ED_270) );
and2 gate( .a(N190), .b(D_54), .O(ED_271) );
and2 gate( .a(N89), .b(D_54_NOT), .O(ED_272) );
and2 gate( .a(N190), .b(D_54), .O(ED_273) );
and2 gate( .a(ED_270), .b(D_55_NOT), .O(ED_274) );
and2 gate( .a(ED_271), .b(D_55), .O(ED_275) );
and2 gate( .a(ED_272), .b(D_55_NOT), .O(ED_276) );
and2 gate( .a(ED_273), .b(D_55), .O(ED_277) );
or2  gate( .a(ED_274), .b(ED_275), .O(ED_278) );
or2  gate( .a(ED_276), .b(ED_278), .O(ED_279) );
or2  gate( .a(ED_279), .b(ED_277), .O(MUX_O_27) );
inv1 gate( .a(D_56),.O(D_56_NOT) );
inv1 gate( .a(D_57),.O(D_57_NOT) );
and2 gate( .a(N14), .b(D_56_NOT), .O(ED_280) );
and2 gate( .a(N420), .b(D_56), .O(ED_281) );
and2 gate( .a(N89), .b(D_56_NOT), .O(ED_282) );
and2 gate( .a(N420), .b(D_56), .O(ED_283) );
and2 gate( .a(ED_280), .b(D_57_NOT), .O(ED_284) );
and2 gate( .a(ED_281), .b(D_57), .O(ED_285) );
and2 gate( .a(ED_282), .b(D_57_NOT), .O(ED_286) );
and2 gate( .a(ED_283), .b(D_57), .O(ED_287) );
or2  gate( .a(ED_284), .b(ED_285), .O(ED_288) );
or2  gate( .a(ED_286), .b(ED_288), .O(ED_289) );
or2  gate( .a(ED_289), .b(ED_287), .O(MUX_O_28) );
inv1 gate( .a(D_58),.O(D_58_NOT) );
inv1 gate( .a(D_59),.O(D_59_NOT) );
and2 gate( .a(N14), .b(D_58_NOT), .O(ED_290) );
and2 gate( .a(N411), .b(D_58), .O(ED_291) );
and2 gate( .a(N89), .b(D_58_NOT), .O(ED_292) );
and2 gate( .a(N411), .b(D_58), .O(ED_293) );
and2 gate( .a(ED_290), .b(D_59_NOT), .O(ED_294) );
and2 gate( .a(ED_291), .b(D_59), .O(ED_295) );
and2 gate( .a(ED_292), .b(D_59_NOT), .O(ED_296) );
and2 gate( .a(ED_293), .b(D_59), .O(ED_297) );
or2  gate( .a(ED_294), .b(ED_295), .O(ED_298) );
or2  gate( .a(ED_296), .b(ED_298), .O(ED_299) );
or2  gate( .a(ED_299), .b(ED_297), .O(MUX_O_29) );
inv1 gate( .a(D_60),.O(D_60_NOT) );
inv1 gate( .a(D_61),.O(D_61_NOT) );
and2 gate( .a(N14), .b(D_60_NOT), .O(ED_300) );
and2 gate( .a(N411), .b(D_60), .O(ED_301) );
and2 gate( .a(N89), .b(D_60_NOT), .O(ED_302) );
and2 gate( .a(N411), .b(D_60), .O(ED_303) );
and2 gate( .a(ED_300), .b(D_61_NOT), .O(ED_304) );
and2 gate( .a(ED_301), .b(D_61), .O(ED_305) );
and2 gate( .a(ED_302), .b(D_61_NOT), .O(ED_306) );
and2 gate( .a(ED_303), .b(D_61), .O(ED_307) );
or2  gate( .a(ED_304), .b(ED_305), .O(ED_308) );
or2  gate( .a(ED_306), .b(ED_308), .O(ED_309) );
or2  gate( .a(ED_309), .b(ED_307), .O(MUX_O_30) );

endmodule