
module c880 (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
             N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
             N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
             N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
             N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
             N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
             N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
             N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
             N865,N866,N874,N878,N879,N880);

input N1_new,N8_new,N13_new,N17_new,N26_new,N29_new,N36_new,N42_new,N51_new,N55_new,
      N59_new,N68_new,N72_new,N73_new,N74_new,N75_new,N80_new,N85_new,N86_new,N87_new,
      N88_new,N89_new,N90_new,N91_new,N96_new,N101_new,N106_new,N111_new,N116_new,N121_new,
      N126_new,N130_new,N135_new,N138_new,N143_new,N146_new,N149_new,N152_new,N153_new,N156_new,
      N159_new,N165_new,N171_new,N177_new,N183_new,N189_new,N195_new,N201_new,N207_new,N210_new,
      N219_new,N228_new,N237_new,N246_new,N255_new,N259_new,N260_new,N261_new,N267_new,N268_new;

input p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,
        p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,
        p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,
        p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,
        p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,
        p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,
        p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,
        p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,
        p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,
        p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,
        p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,
        p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,
        p121,p122,p123,p124,X_1,X_2,X_3,X_4,X_5,X_6,X_7,X_8,X_9,X_10,X_11,X_12,X_13,X_14,X_15,X_16,X_17,X_18,X_19,X_20,X_21,X_22,X_23,X_24,X_25,X_26,X_27,X_28,X_29,X_30,X_31,X_32,X_33,X_34,X_35,X_36,X_37,X_38,X_39,X_40,X_41,X_42,X_43,X_44,X_45,X_46,X_47,X_48,X_49,X_50,X_51,X_52,X_53,X_54,X_55,X_56,X_57,X_58,X_59,X_60,X_61,X_62,X_63,X_64,X_65,X_66,X_67,X_68,X_69,X_70,X_71,X_72,X_73,X_74,X_75,X_76,X_77,X_78,X_79,X_80,X_81,X_82,X_83,X_84,X_85,X_86,X_87,X_88,X_89,X_90,X_91,X_92,X_93,X_94,X_95,X_96,X_97,X_98,X_99,X_100,X_101,X_102,X_103,X_104,X_105,X_106,X_107,X_108,X_109,X_110,X_111,X_112,X_113,X_114,X_115,X_116,X_117,X_118,X_119,X_120,X_121,X_122,X_123,X_124,X_125,X_126,X_127,X_128,X_129,X_130,X_131,X_132,X_133,X_134,X_135,X_136,X_137,X_138,X_139,X_140,X_141,X_142,X_143,X_144,X_145,X_146,X_147,X_148,X_149,X_150,X_151,X_152,X_153,X_154,X_155,X_156,X_157,X_158,X_159,X_160,X_161,X_162,X_163,X_164,X_165,X_166,X_167,X_168,X_169,X_170,X_171,X_172,X_173,X_174,X_175,X_176,X_177,X_178,X_179,X_180,X_181,X_182,X_183,X_184,X_185,X_186,X_187,X_188,X_189,X_190,X_191,X_192,X_193,X_194,X_195,X_196,X_197,X_198,X_199,X_200,X_201,X_202,X_203,X_204,X_205,X_206,X_207,X_208,X_209,X_210,X_211,X_212,X_213,X_214,X_215,X_216,X_217,X_218,X_219,X_220,X_221,X_222,X_223,X_224,X_225,X_226,X_227,X_228,X_229,X_230,X_231,X_232,X_233,X_234,X_235,X_236,X_237,X_238,X_239,X_240,X_241,X_242,X_243,X_244,X_245,X_246,X_247,X_248,X_249,X_250,X_251,X_252,X_253,X_254,X_255,X_256,X_257,X_258,X_259,X_260,X_261,X_262,X_263,X_264,X_265,X_266,X_267,X_268,X_269,X_270,X_271,X_272,X_273,X_274,X_275,X_276,X_277,X_278,X_279,X_280,X_281,X_282,X_283,X_284,X_285,X_286,X_287,X_288;

output N388_new,N389_new,N390_new,N391_new,N418_new,N419_new,N420_new,N421_new,N422_new,N423_new,
       N446_new,N447_new,N448_new,N449_new,N450_new,N767_new,N768_new,N850_new,N863_new,N864_new,
       N865_new,N866_new,N874_new,N878_new,N879_new,N880_new;

wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,
     N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,
     N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,
     N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,
     N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
     N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
     N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,
     N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
     N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
     N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,
     N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,
     N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,
     N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,
     N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
     N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
     N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
     N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,
     N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,
     N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,
     N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,
     N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,
     N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,
     N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,
     N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
     N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
     N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
     N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
     N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,
     N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,
     N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,
     N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,
     N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
     N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
     N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,
     N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,
     N870,N871,N872,N873,N875,N876,N877,
     N101_NOT,N106_NOT,N111_NOT,N116_NOT,N159_NOT,N165_NOT,N171_NOT,N177_NOT,N255_NOT,N259_NOT,
     N280_NOT,N286_NOT,N307_NOT,N308_NOT,N130_NOT,N460_NOT,N130_NOT,N460_NOT,N463_NOT,N135_NOT,
     N91_NOT,N466_NOT,N475_NOT,N476_NOT,N96_NOT,N466_NOT,N451_NOT,N171_NOT,N317_NOT,N506_NOT,
     N510_NOT,N511_NOT,N514_NOT,N515_NOT,N488_NOT,N540_NOT,N246_NOT,N557_NOT,N246_NOT,N569_NOT,
     N587_NOT,N589_NOT,N593_NOT,N590_NOT,N609_NOT,N606_NOT,N228_NOT,N708_NOT,N756_NOT,N732_NOT,
     N700_NOT,N773_NOT,N692_NOT,N796_NOT,N335_NOT,N808_NOT,N682_NOT,N822_NOT,N219_NOT,N842_NOT,
     N417_NOT,N851_NOT,EX1,EX2,EX3,EX4,EX5,EX6,EX7,EX8,EX9,EX10,
     EX11,EX12,EX13,EX14,EX15,EX16,EX17,EX18,EX19,EX20,
     EX21,EX22,EX23,EX24,EX25,EX26,EX27,EX28,EX29,EX30,
     EX31,EX32,EX33,EX34,EX35,EX36,EX37,EX38,EX39,EX40,
     EX41,EX42,EX43,EX44,EX45,EX46,EX47,EX48,EX49,EX50,
     EX51,EX52,EX53,EX54,EX55,EX56,EX57,EX58,EX59,EX60,
     EX61,EX62,EX63,EX64,EX65,EX66,EX67,EX68,EX69,EX70,
     EX71,EX72,EX73,EX74,EX75,EX76,EX77,EX78,EX79,EX80,
     EX81,EX82,EX83,EX84,EX85,EX86,EX87,EX88,EX89,EX90,
     EX91,EX92,EX93,EX94,EX95,EX96,EX97,EX98,EX99,EX100,
     EX101,EX102,EX103,EX104,EX105,EX106,EX107,EX108,EX109,EX110,
     EX111,EX112,EX113,EX114,EX115,EX116,EX117,EX118,EX119,EX120,
     EX121,EX122,EX123,EX124,EX125,EX126,EX127,EX128,EX129,EX130,
     EX131,EX132,EX133,EX134,EX135,EX136,EX137,EX138,EX139,EX140,
     EX141,EX142,EX143,EX144,EX145,EX146,EX147,EX148,EX149,EX150,
     EX151,EX152,EX153,EX154,EX155,EX156,EX157,EX158,EX159,EX160,
     EX161,EX162,EX163,EX164,EX165,EX166,EX167,EX168,EX169,EX170,
     EX171,EX172,EX173,EX174,EX175,EX176,EX177,EX178,EX179,EX180,
     EX181,EX182,EX183,EX184,EX185,EX186,EX187,EX188,EX189,EX190,
     EX191,EX192,EX193,EX194,EX195,EX196,EX197,EX198,EX199,EX200,
     EX201,EX202,EX203,EX204,EX205,EX206,EX207,EX208,EX209,EX210,
     EX211,EX212,EX213,EX214,EX215,EX216,EX217,EX218,EX219,EX220,
     EX221,EX222,EX223,EX224,EX225,EX226,EX227,EX228,EX229,EX230,
     EX231,EX232,EX233,EX234,EX235,EX236,EX237,EX238,EX239,EX240,
     EX241,EX242,EX243,EX244,EX245,EX246,EX247,EX248,EX249,EX250,
     EX251,EX252,EX253,EX254,EX255,EX256,EX257,EX258,EX259,EX260,
     EX261,EX262,EX263,EX264,EX265,EX266,EX267,EX268,EX269,EX270,
     EX271,EX272,EX273,EX274,EX275,EX276,EX277,EX278,EX279,EX280,
     EX281,EX282,EX283,EX284,EX285,EX286,EX287,EX288,EX289,EX290,
     EX291,EX292,EX293,EX294,EX295,EX296,EX297,EX298,EX299,EX300,
     EX301,EX302,EX303,EX304,EX305,EX306,EX307,EX308,EX309,EX310,N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,N865,N866,N874,N878,N879,N880;


nand4 gate1( .a(N1), .b(N8), .c(N13), .d(N17), .O(N269) );
nand4 gate2( .a(N1), .b(N26), .c(N13), .d(N17), .O(N270) );
and3 gate3( .a(N29), .b(N36), .c(N42), .O(N273) );
and3 gate4( .a(N1), .b(N26), .c(N51), .O(N276) );
nand4 gate5( .a(N1), .b(N8), .c(N51), .d(N17), .O(N279) );
nand4 gate6( .a(N1), .b(N8), .c(N13), .d(N55), .O(N280) );
nand4 gate7( .a(N59), .b(N42), .c(N68), .d(N72), .O(N284) );
nand2 gate8( .a(N29), .b(N68), .O(N285) );
nand3 gate9( .a(N59), .b(N68), .c(N74), .O(N286) );
and3 gate10( .a(N29), .b(N75), .c(N80), .O(N287) );
and3 gate11( .a(N29), .b(N75), .c(N42), .O(N290) );
and3 gate12( .a(N29), .b(N36), .c(N80), .O(N291) );
and3 gate13( .a(N29), .b(N36), .c(N42), .O(N292) );
and3 gate14( .a(N59), .b(N75), .c(N80), .O(N293) );
and3 gate15( .a(N59), .b(N75), .c(N42), .O(N294) );
and3 gate16( .a(N59), .b(N36), .c(N80), .O(N295) );
and3 gate17( .a(N59), .b(N36), .c(N42), .O(N296) );
and2 gate18( .a(N85), .b(N86), .O(N297) );
or2 gate19( .a(N87), .b(N88), .O(N298) );
nand2 gate20( .a(N91), .b(N96), .O(N301) );
or2 gate21( .a(N91), .b(N96), .O(N302) );
inv1 gate( .a(N101),.O(N101_NOT) );
inv1 gate( .a(N106),.O(N106_NOT));
and2 gate( .a(N101_NOT), .b(p1), .O(EX1) );
and2 gate( .a(N106_NOT), .b(EX1), .O(EX2) );
and2 gate( .a(N101), .b(p2), .O(EX3) );
and2 gate( .a(N106_NOT), .b(EX3), .O(EX4) );
and2 gate( .a(N101_NOT), .b(p3), .O(EX5) );
and2 gate( .a(N106), .b(EX5), .O(EX6) );
and2 gate( .a(N101), .b(p4), .O(EX7) );
and2 gate( .a(N106), .b(EX7), .O(EX8) );
or2  gate( .a(EX2), .b(EX4), .O(EX9) );
or2  gate( .a(EX6), .b(EX9), .O(EX10) );
or2  gate( .a(EX8), .b(EX10), .O(N303) );
or2 gate23( .a(N101), .b(N106), .O(N304) );
nand2 gate24( .a(N111), .b(N116), .O(N305) );
inv1 gate( .a(N111),.O(N111_NOT) );
inv1 gate( .a(N116),.O(N116_NOT));
and2 gate( .a(N111_NOT), .b(p5), .O(EX11) );
and2 gate( .a(N116_NOT), .b(EX11), .O(EX12) );
and2 gate( .a(N111), .b(p6), .O(EX13) );
and2 gate( .a(N116_NOT), .b(EX13), .O(EX14) );
and2 gate( .a(N111_NOT), .b(p7), .O(EX15) );
and2 gate( .a(N116), .b(EX15), .O(EX16) );
and2 gate( .a(N111), .b(p8), .O(EX17) );
and2 gate( .a(N116), .b(EX17), .O(EX18) );
or2  gate( .a(EX12), .b(EX14), .O(EX19) );
or2  gate( .a(EX16), .b(EX19), .O(EX20) );
or2  gate( .a(EX18), .b(EX20), .O(N306) );
nand2 gate26( .a(N121), .b(N126), .O(N307) );
or2 gate27( .a(N121), .b(N126), .O(N308) );
and2 gate28( .a(N8), .b(N138), .O(N309) );
inv1 gate29( .a(N268), .O(N310) );
and2 gate30( .a(N51), .b(N138), .O(N316) );
and2 gate31( .a(N17), .b(N138), .O(N317) );
and2 gate32( .a(N152), .b(N138), .O(N318) );
nand2 gate33( .a(N59), .b(N156), .O(N319) );
nor2 gate34( .a(N17), .b(N42), .O(N322) );
and2 gate35( .a(N17), .b(N42), .O(N323) );
nand2 gate36( .a(N159), .b(N165), .O(N324) );
inv1 gate( .a(N159),.O(N159_NOT) );
inv1 gate( .a(N165),.O(N165_NOT));
and2 gate( .a(N159_NOT), .b(p9), .O(EX21) );
and2 gate( .a(N165_NOT), .b(EX21), .O(EX22) );
and2 gate( .a(N159), .b(p10), .O(EX23) );
and2 gate( .a(N165_NOT), .b(EX23), .O(EX24) );
and2 gate( .a(N159_NOT), .b(p11), .O(EX25) );
and2 gate( .a(N165), .b(EX25), .O(EX26) );
and2 gate( .a(N159), .b(p12), .O(EX27) );
and2 gate( .a(N165), .b(EX27), .O(EX28) );
or2  gate( .a(EX22), .b(EX24), .O(EX29) );
or2  gate( .a(EX26), .b(EX29), .O(EX30) );
or2  gate( .a(EX28), .b(EX30), .O(N325) );
inv1 gate( .a(N171),.O(N171_NOT) );
inv1 gate( .a(N177),.O(N177_NOT));
and2 gate( .a(N171_NOT), .b(p13), .O(EX31) );
and2 gate( .a(N177_NOT), .b(EX31), .O(EX32) );
and2 gate( .a(N171), .b(p14), .O(EX33) );
and2 gate( .a(N177_NOT), .b(EX33), .O(EX34) );
and2 gate( .a(N171_NOT), .b(p15), .O(EX35) );
and2 gate( .a(N177), .b(EX35), .O(EX36) );
and2 gate( .a(N171), .b(p16), .O(EX37) );
and2 gate( .a(N177), .b(EX37), .O(EX38) );
or2  gate( .a(EX32), .b(EX34), .O(EX39) );
or2  gate( .a(EX36), .b(EX39), .O(EX40) );
or2  gate( .a(EX38), .b(EX40), .O(N326) );
or2 gate39( .a(N171), .b(N177), .O(N327) );
nand2 gate40( .a(N183), .b(N189), .O(N328) );
or2 gate41( .a(N183), .b(N189), .O(N329) );
nand2 gate42( .a(N195), .b(N201), .O(N330) );
or2 gate43( .a(N195), .b(N201), .O(N331) );
and2 gate44( .a(N210), .b(N91), .O(N332) );
and2 gate45( .a(N210), .b(N96), .O(N333) );
and2 gate46( .a(N210), .b(N101), .O(N334) );
and2 gate47( .a(N210), .b(N106), .O(N335) );
and2 gate48( .a(N210), .b(N111), .O(N336) );
inv1 gate( .a(N255),.O(N255_NOT) );
inv1 gate( .a(N259),.O(N259_NOT));
and2 gate( .a(N255_NOT), .b(p17), .O(EX41) );
and2 gate( .a(N259_NOT), .b(EX41), .O(EX42) );
and2 gate( .a(N255), .b(p18), .O(EX43) );
and2 gate( .a(N259_NOT), .b(EX43), .O(EX44) );
and2 gate( .a(N255_NOT), .b(p19), .O(EX45) );
and2 gate( .a(N259), .b(EX45), .O(EX46) );
and2 gate( .a(N255), .b(p20), .O(EX47) );
and2 gate( .a(N259), .b(EX47), .O(EX48) );
or2  gate( .a(EX42), .b(EX44), .O(EX49) );
or2  gate( .a(EX46), .b(EX49), .O(EX50) );
or2  gate( .a(EX48), .b(EX50), .O(N337) );
and2 gate50( .a(N210), .b(N116), .O(N338) );
and2 gate51( .a(N255), .b(N260), .O(N339) );
and2 gate52( .a(N210), .b(N121), .O(N340) );
and2 gate53( .a(N255), .b(N267), .O(N341) );
inv1 gate54( .a(N269), .O(N342) );
inv1 gate55( .a(N273), .O(N343) );
or2 gate56( .a(N270), .b(N273), .O(N344) );
inv1 gate57( .a(N276), .O(N345) );
inv1 gate58( .a(N276), .O(N346) );
inv1 gate59( .a(N279), .O(N347) );
nor2 gate60( .a(N280), .b(N284), .O(N348) );
or2 gate61( .a(N280), .b(N285), .O(N349) );
inv1 gate( .a(N280),.O(N280_NOT) );
inv1 gate( .a(N286),.O(N286_NOT));
and2 gate( .a(N280_NOT), .b(p21), .O(EX51) );
and2 gate( .a(N286_NOT), .b(EX51), .O(EX52) );
and2 gate( .a(N280), .b(p22), .O(EX53) );
and2 gate( .a(N286_NOT), .b(EX53), .O(EX54) );
and2 gate( .a(N280_NOT), .b(p23), .O(EX55) );
and2 gate( .a(N286), .b(EX55), .O(EX56) );
and2 gate( .a(N280), .b(p24), .O(EX57) );
and2 gate( .a(N286), .b(EX57), .O(EX58) );
or2  gate( .a(EX52), .b(EX54), .O(EX59) );
or2  gate( .a(EX56), .b(EX59), .O(EX60) );
or2  gate( .a(EX58), .b(EX60), .O(N350) );
inv1 gate63( .a(N293), .O(N351) );
inv1 gate64( .a(N294), .O(N352) );
inv1 gate65( .a(N295), .O(N353) );
inv1 gate66( .a(N296), .O(N354) );
nand2 gate67( .a(N89), .b(N298), .O(N355) );
and2 gate68( .a(N90), .b(N298), .O(N356) );
nand2 gate69( .a(N301), .b(N302), .O(N357) );
nand2 gate70( .a(N303), .b(N304), .O(N360) );
nand2 gate71( .a(N305), .b(N306), .O(N363) );
inv1 gate( .a(N307),.O(N307_NOT) );
inv1 gate( .a(N308),.O(N308_NOT));
and2 gate( .a(N307_NOT), .b(p25), .O(EX61) );
and2 gate( .a(N308_NOT), .b(EX61), .O(EX62) );
and2 gate( .a(N307), .b(p26), .O(EX63) );
and2 gate( .a(N308_NOT), .b(EX63), .O(EX64) );
and2 gate( .a(N307_NOT), .b(p27), .O(EX65) );
and2 gate( .a(N308), .b(EX65), .O(EX66) );
and2 gate( .a(N307), .b(p28), .O(EX67) );
and2 gate( .a(N308), .b(EX67), .O(EX68) );
or2  gate( .a(EX62), .b(EX64), .O(EX69) );
or2  gate( .a(EX66), .b(EX69), .O(EX70) );
or2  gate( .a(EX68), .b(EX70), .O(N366) );
inv1 gate73( .a(N310), .O(N369) );
nor2 gate74( .a(N322), .b(N323), .O(N375) );
nand2 gate75( .a(N324), .b(N325), .O(N376) );
nand2 gate76( .a(N326), .b(N327), .O(N379) );
nand2 gate77( .a(N328), .b(N329), .O(N382) );
nand2 gate78( .a(N330), .b(N331), .O(N385) );
buf1 gate79( .a(N290), .O(N388) );
buf1 gate80( .a(N291), .O(N389) );
buf1 gate81( .a(N292), .O(N390) );
buf1 gate82( .a(N297), .O(N391) );
or2 gate83( .a(N270), .b(N343), .O(N392) );
inv1 gate84( .a(N345), .O(N393) );
inv1 gate85( .a(N346), .O(N399) );
and2 gate86( .a(N348), .b(N73), .O(N400) );
inv1 gate87( .a(N349), .O(N401) );
inv1 gate88( .a(N350), .O(N402) );
inv1 gate89( .a(N355), .O(N403) );
inv1 gate90( .a(N357), .O(N404) );
inv1 gate91( .a(N360), .O(N405) );
and2 gate92( .a(N357), .b(N360), .O(N406) );
inv1 gate93( .a(N363), .O(N407) );
inv1 gate94( .a(N366), .O(N408) );
and2 gate95( .a(N363), .b(N366), .O(N409) );
nand2 gate96( .a(N347), .b(N352), .O(N410) );
inv1 gate97( .a(N376), .O(N411) );
inv1 gate98( .a(N379), .O(N412) );
and2 gate99( .a(N376), .b(N379), .O(N413) );
inv1 gate100( .a(N382), .O(N414) );
inv1 gate101( .a(N385), .O(N415) );
and2 gate102( .a(N382), .b(N385), .O(N416) );
and2 gate103( .a(N210), .b(N369), .O(N417) );
buf1 gate104( .a(N342), .O(N418) );
buf1 gate105( .a(N344), .O(N419) );
buf1 gate106( .a(N351), .O(N420) );
buf1 gate107( .a(N353), .O(N421) );
buf1 gate108( .a(N354), .O(N422) );
buf1 gate109( .a(N356), .O(N423) );
inv1 gate110( .a(N400), .O(N424) );
and2 gate111( .a(N404), .b(N405), .O(N425) );
and2 gate112( .a(N407), .b(N408), .O(N426) );
and3 gate113( .a(N319), .b(N393), .c(N55), .O(N427) );
and3 gate114( .a(N393), .b(N17), .c(N287), .O(N432) );
nand3 gate115( .a(N393), .b(N287), .c(N55), .O(N437) );
nand4 gate116( .a(N375), .b(N59), .c(N156), .d(N393), .O(N442) );
nand3 gate117( .a(N393), .b(N319), .c(N17), .O(N443) );
and2 gate118( .a(N411), .b(N412), .O(N444) );
and2 gate119( .a(N414), .b(N415), .O(N445) );
buf1 gate120( .a(N392), .O(N446) );
buf1 gate121( .a(N399), .O(N447) );
buf1 gate122( .a(N401), .O(N448) );
buf1 gate123( .a(N402), .O(N449) );
buf1 gate124( .a(N403), .O(N450) );
inv1 gate125( .a(N424), .O(N451) );
nor2 gate126( .a(N406), .b(N425), .O(N460) );
nor2 gate127( .a(N409), .b(N426), .O(N463) );
nand2 gate128( .a(N442), .b(N410), .O(N466) );
and2 gate129( .a(N143), .b(N427), .O(N475) );
and2 gate130( .a(N310), .b(N432), .O(N476) );
and2 gate131( .a(N146), .b(N427), .O(N477) );
and2 gate132( .a(N310), .b(N432), .O(N478) );
and2 gate133( .a(N149), .b(N427), .O(N479) );
and2 gate134( .a(N310), .b(N432), .O(N480) );
and2 gate135( .a(N153), .b(N427), .O(N481) );
and2 gate136( .a(N310), .b(N432), .O(N482) );
nand2 gate137( .a(N443), .b(N1), .O(N483) );
or2 gate138( .a(N369), .b(N437), .O(N488) );
or2 gate139( .a(N369), .b(N437), .O(N489) );
or2 gate140( .a(N369), .b(N437), .O(N490) );
or2 gate141( .a(N369), .b(N437), .O(N491) );
nor2 gate142( .a(N413), .b(N444), .O(N492) );
nor2 gate143( .a(N416), .b(N445), .O(N495) );
inv1 gate( .a(N130),.O(N130_NOT) );
inv1 gate( .a(N460),.O(N460_NOT));
and2 gate( .a(N130_NOT), .b(p29), .O(EX71) );
and2 gate( .a(N460_NOT), .b(EX71), .O(EX72) );
and2 gate( .a(N130), .b(p30), .O(EX73) );
and2 gate( .a(N460_NOT), .b(EX73), .O(EX74) );
and2 gate( .a(N130_NOT), .b(p31), .O(EX75) );
and2 gate( .a(N460), .b(EX75), .O(EX76) );
and2 gate( .a(N130), .b(p32), .O(EX77) );
and2 gate( .a(N460), .b(EX77), .O(EX78) );
or2  gate( .a(EX72), .b(EX74), .O(EX79) );
or2  gate( .a(EX76), .b(EX79), .O(EX80) );
or2  gate( .a(EX78), .b(EX80), .O(N498) );
inv1 gate( .a(N130),.O(N130_NOT) );
inv1 gate( .a(N460),.O(N460_NOT));
and2 gate( .a(N130_NOT), .b(p33), .O(EX81) );
and2 gate( .a(N460_NOT), .b(EX81), .O(EX82) );
and2 gate( .a(N130), .b(p34), .O(EX83) );
and2 gate( .a(N460_NOT), .b(EX83), .O(EX84) );
and2 gate( .a(N130_NOT), .b(p35), .O(EX85) );
and2 gate( .a(N460), .b(EX85), .O(EX86) );
and2 gate( .a(N130), .b(p36), .O(EX87) );
and2 gate( .a(N460), .b(EX87), .O(EX88) );
or2  gate( .a(EX82), .b(EX84), .O(EX89) );
or2  gate( .a(EX86), .b(EX89), .O(EX90) );
or2  gate( .a(EX88), .b(EX90), .O(N499) );
inv1 gate( .a(N463),.O(N463_NOT) );
inv1 gate( .a(N135),.O(N135_NOT));
and2 gate( .a(N463_NOT), .b(p37), .O(EX91) );
and2 gate( .a(N135_NOT), .b(EX91), .O(EX92) );
and2 gate( .a(N463), .b(p38), .O(EX93) );
and2 gate( .a(N135_NOT), .b(EX93), .O(EX94) );
and2 gate( .a(N463_NOT), .b(p39), .O(EX95) );
and2 gate( .a(N135), .b(EX95), .O(EX96) );
and2 gate( .a(N463), .b(p40), .O(EX97) );
and2 gate( .a(N135), .b(EX97), .O(EX98) );
or2  gate( .a(EX92), .b(EX94), .O(EX99) );
or2  gate( .a(EX96), .b(EX99), .O(EX100) );
or2  gate( .a(EX98), .b(EX100), .O(N500) );
or2 gate147( .a(N463), .b(N135), .O(N501) );
inv1 gate( .a(N91),.O(N91_NOT) );
inv1 gate( .a(N466),.O(N466_NOT));
and2 gate( .a(N91_NOT), .b(p41), .O(EX101) );
and2 gate( .a(N466_NOT), .b(EX101), .O(EX102) );
and2 gate( .a(N91), .b(p42), .O(EX103) );
and2 gate( .a(N466_NOT), .b(EX103), .O(EX104) );
and2 gate( .a(N91_NOT), .b(p43), .O(EX105) );
and2 gate( .a(N466), .b(EX105), .O(EX106) );
and2 gate( .a(N91), .b(p44), .O(EX107) );
and2 gate( .a(N466), .b(EX107), .O(EX108) );
or2  gate( .a(EX102), .b(EX104), .O(EX109) );
or2  gate( .a(EX106), .b(EX109), .O(EX110) );
or2  gate( .a(EX108), .b(EX110), .O(N502) );
inv1 gate( .a(N475),.O(N475_NOT) );
inv1 gate( .a(N476),.O(N476_NOT));
and2 gate( .a(N475_NOT), .b(p45), .O(EX111) );
and2 gate( .a(N476_NOT), .b(EX111), .O(EX112) );
and2 gate( .a(N475), .b(p46), .O(EX113) );
and2 gate( .a(N476_NOT), .b(EX113), .O(EX114) );
and2 gate( .a(N475_NOT), .b(p47), .O(EX115) );
and2 gate( .a(N476), .b(EX115), .O(EX116) );
and2 gate( .a(N475), .b(p48), .O(EX117) );
and2 gate( .a(N476), .b(EX117), .O(EX118) );
or2  gate( .a(EX112), .b(EX114), .O(EX119) );
or2  gate( .a(EX116), .b(EX119), .O(EX120) );
or2  gate( .a(EX118), .b(EX120), .O(N503) );
inv1 gate( .a(N96),.O(N96_NOT) );
inv1 gate( .a(N466),.O(N466_NOT));
and2 gate( .a(N96_NOT), .b(p49), .O(EX121) );
and2 gate( .a(N466_NOT), .b(EX121), .O(EX122) );
and2 gate( .a(N96), .b(p50), .O(EX123) );
and2 gate( .a(N466_NOT), .b(EX123), .O(EX124) );
and2 gate( .a(N96_NOT), .b(p51), .O(EX125) );
and2 gate( .a(N466), .b(EX125), .O(EX126) );
and2 gate( .a(N96), .b(p52), .O(EX127) );
and2 gate( .a(N466), .b(EX127), .O(EX128) );
or2  gate( .a(EX122), .b(EX124), .O(EX129) );
or2  gate( .a(EX126), .b(EX129), .O(EX130) );
or2  gate( .a(EX128), .b(EX130), .O(N504) );
nor2 gate151( .a(N477), .b(N478), .O(N505) );
and2 gate152( .a(N101), .b(N466), .O(N506) );
nor2 gate153( .a(N479), .b(N480), .O(N507) );
and2 gate154( .a(N106), .b(N466), .O(N508) );
nor2 gate155( .a(N481), .b(N482), .O(N509) );
and2 gate156( .a(N143), .b(N483), .O(N510) );
and2 gate157( .a(N111), .b(N466), .O(N511) );
and2 gate158( .a(N146), .b(N483), .O(N512) );
and2 gate159( .a(N116), .b(N466), .O(N513) );
and2 gate160( .a(N149), .b(N483), .O(N514) );
and2 gate161( .a(N121), .b(N466), .O(N515) );
and2 gate162( .a(N153), .b(N483), .O(N516) );
and2 gate163( .a(N126), .b(N466), .O(N517) );
nand2 gate164( .a(N130), .b(N492), .O(N518) );
or2 gate165( .a(N130), .b(N492), .O(N519) );
nand2 gate166( .a(N495), .b(N207), .O(N520) );
or2 gate167( .a(N495), .b(N207), .O(N521) );
and2 gate168( .a(N451), .b(N159), .O(N522) );
and2 gate169( .a(N451), .b(N165), .O(N523) );
inv1 gate( .a(N451),.O(N451_NOT) );
inv1 gate( .a(N171),.O(N171_NOT));
and2 gate( .a(N451_NOT), .b(p53), .O(EX131) );
and2 gate( .a(N171_NOT), .b(EX131), .O(EX132) );
and2 gate( .a(N451), .b(p54), .O(EX133) );
and2 gate( .a(N171_NOT), .b(EX133), .O(EX134) );
and2 gate( .a(N451_NOT), .b(p55), .O(EX135) );
and2 gate( .a(N171), .b(EX135), .O(EX136) );
and2 gate( .a(N451), .b(p56), .O(EX137) );
and2 gate( .a(N171), .b(EX137), .O(EX138) );
or2  gate( .a(EX132), .b(EX134), .O(EX139) );
or2  gate( .a(EX136), .b(EX139), .O(EX140) );
or2  gate( .a(EX138), .b(EX140), .O(N524) );
and2 gate171( .a(N451), .b(N177), .O(N525) );
and2 gate172( .a(N451), .b(N183), .O(N526) );
nand2 gate173( .a(N451), .b(N189), .O(N527) );
nand2 gate174( .a(N451), .b(N195), .O(N528) );
nand2 gate175( .a(N451), .b(N201), .O(N529) );
nand2 gate176( .a(N498), .b(N499), .O(N530) );
nand2 gate177( .a(N500), .b(N501), .O(N533) );
nor2 gate178( .a(N309), .b(N502), .O(N536) );
nor2 gate179( .a(N316), .b(N504), .O(N537) );
inv1 gate( .a(N317),.O(N317_NOT) );
inv1 gate( .a(N506),.O(N506_NOT));
and2 gate( .a(N317_NOT), .b(p57), .O(EX141) );
and2 gate( .a(N506_NOT), .b(EX141), .O(EX142) );
and2 gate( .a(N317), .b(p58), .O(EX143) );
and2 gate( .a(N506_NOT), .b(EX143), .O(EX144) );
and2 gate( .a(N317_NOT), .b(p59), .O(EX145) );
and2 gate( .a(N506), .b(EX145), .O(EX146) );
and2 gate( .a(N317), .b(p60), .O(EX147) );
and2 gate( .a(N506), .b(EX147), .O(EX148) );
or2  gate( .a(EX142), .b(EX144), .O(EX149) );
or2  gate( .a(EX146), .b(EX149), .O(EX150) );
or2  gate( .a(EX148), .b(EX150), .O(N538) );
nor2 gate181( .a(N318), .b(N508), .O(N539) );
inv1 gate( .a(N510),.O(N510_NOT) );
inv1 gate( .a(N511),.O(N511_NOT));
and2 gate( .a(N510_NOT), .b(p61), .O(EX151) );
and2 gate( .a(N511_NOT), .b(EX151), .O(EX152) );
and2 gate( .a(N510), .b(p62), .O(EX153) );
and2 gate( .a(N511_NOT), .b(EX153), .O(EX154) );
and2 gate( .a(N510_NOT), .b(p63), .O(EX155) );
and2 gate( .a(N511), .b(EX155), .O(EX156) );
and2 gate( .a(N510), .b(p64), .O(EX157) );
and2 gate( .a(N511), .b(EX157), .O(EX158) );
or2  gate( .a(EX152), .b(EX154), .O(EX159) );
or2  gate( .a(EX156), .b(EX159), .O(EX160) );
or2  gate( .a(EX158), .b(EX160), .O(N540) );
nor2 gate183( .a(N512), .b(N513), .O(N541) );
inv1 gate( .a(N514),.O(N514_NOT) );
inv1 gate( .a(N515),.O(N515_NOT));
and2 gate( .a(N514_NOT), .b(p65), .O(EX161) );
and2 gate( .a(N515_NOT), .b(EX161), .O(EX162) );
and2 gate( .a(N514), .b(p66), .O(EX163) );
and2 gate( .a(N515_NOT), .b(EX163), .O(EX164) );
and2 gate( .a(N514_NOT), .b(p67), .O(EX165) );
and2 gate( .a(N515), .b(EX165), .O(EX166) );
and2 gate( .a(N514), .b(p68), .O(EX167) );
and2 gate( .a(N515), .b(EX167), .O(EX168) );
or2  gate( .a(EX162), .b(EX164), .O(EX169) );
or2  gate( .a(EX166), .b(EX169), .O(EX170) );
or2  gate( .a(EX168), .b(EX170), .O(N542) );
nor2 gate185( .a(N516), .b(N517), .O(N543) );
nand2 gate186( .a(N518), .b(N519), .O(N544) );
nand2 gate187( .a(N520), .b(N521), .O(N547) );
inv1 gate188( .a(N530), .O(N550) );
inv1 gate189( .a(N533), .O(N551) );
and2 gate190( .a(N530), .b(N533), .O(N552) );
nand2 gate191( .a(N536), .b(N503), .O(N553) );
nand2 gate192( .a(N537), .b(N505), .O(N557) );
nand2 gate193( .a(N538), .b(N507), .O(N561) );
nand2 gate194( .a(N539), .b(N509), .O(N565) );
inv1 gate( .a(N488),.O(N488_NOT) );
inv1 gate( .a(N540),.O(N540_NOT));
and2 gate( .a(N488_NOT), .b(p69), .O(EX171) );
and2 gate( .a(N540_NOT), .b(EX171), .O(EX172) );
and2 gate( .a(N488), .b(p70), .O(EX173) );
and2 gate( .a(N540_NOT), .b(EX173), .O(EX174) );
and2 gate( .a(N488_NOT), .b(p71), .O(EX175) );
and2 gate( .a(N540), .b(EX175), .O(EX176) );
and2 gate( .a(N488), .b(p72), .O(EX177) );
and2 gate( .a(N540), .b(EX177), .O(EX178) );
or2  gate( .a(EX172), .b(EX174), .O(EX179) );
or2  gate( .a(EX176), .b(EX179), .O(EX180) );
or2  gate( .a(EX178), .b(EX180), .O(N569) );
nand2 gate196( .a(N489), .b(N541), .O(N573) );
nand2 gate197( .a(N490), .b(N542), .O(N577) );
nand2 gate198( .a(N491), .b(N543), .O(N581) );
inv1 gate199( .a(N544), .O(N585) );
inv1 gate200( .a(N547), .O(N586) );
and2 gate201( .a(N544), .b(N547), .O(N587) );
and2 gate202( .a(N550), .b(N551), .O(N588) );
and2 gate203( .a(N585), .b(N586), .O(N589) );
nand2 gate204( .a(N553), .b(N159), .O(N590) );
or2 gate205( .a(N553), .b(N159), .O(N593) );
and2 gate206( .a(N246), .b(N553), .O(N596) );
nand2 gate207( .a(N557), .b(N165), .O(N597) );
or2 gate208( .a(N557), .b(N165), .O(N600) );
inv1 gate( .a(N246),.O(N246_NOT) );
inv1 gate( .a(N557),.O(N557_NOT));
and2 gate( .a(N246_NOT), .b(p73), .O(EX181) );
and2 gate( .a(N557_NOT), .b(EX181), .O(EX182) );
and2 gate( .a(N246), .b(p74), .O(EX183) );
and2 gate( .a(N557_NOT), .b(EX183), .O(EX184) );
and2 gate( .a(N246_NOT), .b(p75), .O(EX185) );
and2 gate( .a(N557), .b(EX185), .O(EX186) );
and2 gate( .a(N246), .b(p76), .O(EX187) );
and2 gate( .a(N557), .b(EX187), .O(EX188) );
or2  gate( .a(EX182), .b(EX184), .O(EX189) );
or2  gate( .a(EX186), .b(EX189), .O(EX190) );
or2  gate( .a(EX188), .b(EX190), .O(N605) );
nand2 gate210( .a(N561), .b(N171), .O(N606) );
or2 gate211( .a(N561), .b(N171), .O(N609) );
and2 gate212( .a(N246), .b(N561), .O(N615) );
nand2 gate213( .a(N565), .b(N177), .O(N616) );
or2 gate214( .a(N565), .b(N177), .O(N619) );
and2 gate215( .a(N246), .b(N565), .O(N624) );
nand2 gate216( .a(N569), .b(N183), .O(N625) );
or2 gate217( .a(N569), .b(N183), .O(N628) );
inv1 gate( .a(N246),.O(N246_NOT) );
inv1 gate( .a(N569),.O(N569_NOT));
and2 gate( .a(N246_NOT), .b(p77), .O(EX191) );
and2 gate( .a(N569_NOT), .b(EX191), .O(EX192) );
and2 gate( .a(N246), .b(p78), .O(EX193) );
and2 gate( .a(N569_NOT), .b(EX193), .O(EX194) );
and2 gate( .a(N246_NOT), .b(p79), .O(EX195) );
and2 gate( .a(N569), .b(EX195), .O(EX196) );
and2 gate( .a(N246), .b(p80), .O(EX197) );
and2 gate( .a(N569), .b(EX197), .O(EX198) );
or2  gate( .a(EX192), .b(EX194), .O(EX199) );
or2  gate( .a(EX196), .b(EX199), .O(EX200) );
or2  gate( .a(EX198), .b(EX200), .O(N631) );
nand2 gate219( .a(N573), .b(N189), .O(N632) );
or2 gate220( .a(N573), .b(N189), .O(N635) );
and2 gate221( .a(N246), .b(N573), .O(N640) );
nand2 gate222( .a(N577), .b(N195), .O(N641) );
or2 gate223( .a(N577), .b(N195), .O(N644) );
and2 gate224( .a(N246), .b(N577), .O(N650) );
nand2 gate225( .a(N581), .b(N201), .O(N651) );
or2 gate226( .a(N581), .b(N201), .O(N654) );
and2 gate227( .a(N246), .b(N581), .O(N659) );
nor2 gate228( .a(N552), .b(N588), .O(N660) );
inv1 gate( .a(N587),.O(N587_NOT) );
inv1 gate( .a(N589),.O(N589_NOT));
and2 gate( .a(N587_NOT), .b(p81), .O(EX201) );
and2 gate( .a(N589_NOT), .b(EX201), .O(EX202) );
and2 gate( .a(N587), .b(p82), .O(EX203) );
and2 gate( .a(N589_NOT), .b(EX203), .O(EX204) );
and2 gate( .a(N587_NOT), .b(p83), .O(EX205) );
and2 gate( .a(N589), .b(EX205), .O(EX206) );
and2 gate( .a(N587), .b(p84), .O(EX207) );
and2 gate( .a(N589), .b(EX207), .O(EX208) );
or2  gate( .a(EX202), .b(EX204), .O(EX209) );
or2  gate( .a(EX206), .b(EX209), .O(EX210) );
or2  gate( .a(EX208), .b(EX210), .O(N661) );
inv1 gate230( .a(N590), .O(N662) );
inv1 gate( .a(N593),.O(N593_NOT) );
inv1 gate( .a(N590),.O(N590_NOT));
and2 gate( .a(N593_NOT), .b(p85), .O(EX211) );
and2 gate( .a(N590_NOT), .b(EX211), .O(EX212) );
and2 gate( .a(N593), .b(p86), .O(EX213) );
and2 gate( .a(N590_NOT), .b(EX213), .O(EX214) );
and2 gate( .a(N593_NOT), .b(p87), .O(EX215) );
and2 gate( .a(N590), .b(EX215), .O(EX216) );
and2 gate( .a(N593), .b(p88), .O(EX217) );
and2 gate( .a(N590), .b(EX217), .O(EX218) );
or2  gate( .a(EX212), .b(EX214), .O(EX219) );
or2  gate( .a(EX216), .b(EX219), .O(EX220) );
or2  gate( .a(EX218), .b(EX220), .O(N665) );
nor2 gate232( .a(N596), .b(N522), .O(N669) );
inv1 gate233( .a(N597), .O(N670) );
and2 gate234( .a(N600), .b(N597), .O(N673) );
nor2 gate235( .a(N605), .b(N523), .O(N677) );
inv1 gate236( .a(N606), .O(N678) );
inv1 gate( .a(N609),.O(N609_NOT) );
inv1 gate( .a(N606),.O(N606_NOT));
and2 gate( .a(N609_NOT), .b(p89), .O(EX221) );
and2 gate( .a(N606_NOT), .b(EX221), .O(EX222) );
and2 gate( .a(N609), .b(p90), .O(EX223) );
and2 gate( .a(N606_NOT), .b(EX223), .O(EX224) );
and2 gate( .a(N609_NOT), .b(p91), .O(EX225) );
and2 gate( .a(N606), .b(EX225), .O(EX226) );
and2 gate( .a(N609), .b(p92), .O(EX227) );
and2 gate( .a(N606), .b(EX227), .O(EX228) );
or2  gate( .a(EX222), .b(EX224), .O(EX229) );
or2  gate( .a(EX226), .b(EX229), .O(EX230) );
or2  gate( .a(EX228), .b(EX230), .O(N682) );
nor2 gate238( .a(N615), .b(N524), .O(N686) );
inv1 gate239( .a(N616), .O(N687) );
and2 gate240( .a(N619), .b(N616), .O(N692) );
nor2 gate241( .a(N624), .b(N525), .O(N696) );
inv1 gate242( .a(N625), .O(N697) );
and2 gate243( .a(N628), .b(N625), .O(N700) );
nor2 gate244( .a(N631), .b(N526), .O(N704) );
inv1 gate245( .a(N632), .O(N705) );
and2 gate246( .a(N635), .b(N632), .O(N708) );
nor2 gate247( .a(N337), .b(N640), .O(N712) );
inv1 gate248( .a(N641), .O(N713) );
and2 gate249( .a(N644), .b(N641), .O(N717) );
nor2 gate250( .a(N339), .b(N650), .O(N721) );
inv1 gate251( .a(N651), .O(N722) );
and2 gate252( .a(N654), .b(N651), .O(N727) );
nor2 gate253( .a(N341), .b(N659), .O(N731) );
nand2 gate254( .a(N654), .b(N261), .O(N732) );
nand3 gate255( .a(N644), .b(N654), .c(N261), .O(N733) );
nand4 gate256( .a(N635), .b(N644), .c(N654), .d(N261), .O(N734) );
inv1 gate257( .a(N662), .O(N735) );
and2 gate258( .a(N228), .b(N665), .O(N736) );
and2 gate259( .a(N237), .b(N662), .O(N737) );
inv1 gate260( .a(N670), .O(N738) );
and2 gate261( .a(N228), .b(N673), .O(N739) );
and2 gate262( .a(N237), .b(N670), .O(N740) );
inv1 gate263( .a(N678), .O(N741) );
and2 gate264( .a(N228), .b(N682), .O(N742) );
and2 gate265( .a(N237), .b(N678), .O(N743) );
inv1 gate266( .a(N687), .O(N744) );
and2 gate267( .a(N228), .b(N692), .O(N745) );
and2 gate268( .a(N237), .b(N687), .O(N746) );
inv1 gate269( .a(N697), .O(N747) );
and2 gate270( .a(N228), .b(N700), .O(N748) );
and2 gate271( .a(N237), .b(N697), .O(N749) );
inv1 gate272( .a(N705), .O(N750) );
inv1 gate( .a(N228),.O(N228_NOT) );
inv1 gate( .a(N708),.O(N708_NOT));
and2 gate( .a(N228_NOT), .b(p93), .O(EX231) );
and2 gate( .a(N708_NOT), .b(EX231), .O(EX232) );
and2 gate( .a(N228), .b(p94), .O(EX233) );
and2 gate( .a(N708_NOT), .b(EX233), .O(EX234) );
and2 gate( .a(N228_NOT), .b(p95), .O(EX235) );
and2 gate( .a(N708), .b(EX235), .O(EX236) );
and2 gate( .a(N228), .b(p96), .O(EX237) );
and2 gate( .a(N708), .b(EX237), .O(EX238) );
or2  gate( .a(EX232), .b(EX234), .O(EX239) );
or2  gate( .a(EX236), .b(EX239), .O(EX240) );
or2  gate( .a(EX238), .b(EX240), .O(N751) );
and2 gate274( .a(N237), .b(N705), .O(N752) );
inv1 gate275( .a(N713), .O(N753) );
and2 gate276( .a(N228), .b(N717), .O(N754) );
and2 gate277( .a(N237), .b(N713), .O(N755) );
inv1 gate278( .a(N722), .O(N756) );
nor2 gate279( .a(N727), .b(N261), .O(N757) );
and2 gate280( .a(N727), .b(N261), .O(N758) );
and2 gate281( .a(N228), .b(N727), .O(N759) );
and2 gate282( .a(N237), .b(N722), .O(N760) );
nand2 gate283( .a(N644), .b(N722), .O(N761) );
nand2 gate284( .a(N635), .b(N713), .O(N762) );
nand3 gate285( .a(N635), .b(N644), .c(N722), .O(N763) );
nand2 gate286( .a(N609), .b(N687), .O(N764) );
nand2 gate287( .a(N600), .b(N678), .O(N765) );
nand3 gate288( .a(N600), .b(N609), .c(N687), .O(N766) );
buf1 gate289( .a(N660), .O(N767) );
buf1 gate290( .a(N661), .O(N768) );
nor2 gate291( .a(N736), .b(N737), .O(N769) );
nor2 gate292( .a(N739), .b(N740), .O(N770) );
nor2 gate293( .a(N742), .b(N743), .O(N771) );
nor2 gate294( .a(N745), .b(N746), .O(N772) );
nand4 gate295( .a(N750), .b(N762), .c(N763), .d(N734), .O(N773) );
nor2 gate296( .a(N748), .b(N749), .O(N777) );
nand3 gate297( .a(N753), .b(N761), .c(N733), .O(N778) );
nor2 gate298( .a(N751), .b(N752), .O(N781) );
inv1 gate( .a(N756),.O(N756_NOT) );
inv1 gate( .a(N732),.O(N732_NOT));
and2 gate( .a(N756_NOT), .b(p97), .O(EX241) );
and2 gate( .a(N732_NOT), .b(EX241), .O(EX242) );
and2 gate( .a(N756), .b(p98), .O(EX243) );
and2 gate( .a(N732_NOT), .b(EX243), .O(EX244) );
and2 gate( .a(N756_NOT), .b(p99), .O(EX245) );
and2 gate( .a(N732), .b(EX245), .O(EX246) );
and2 gate( .a(N756), .b(p100), .O(EX247) );
and2 gate( .a(N732), .b(EX247), .O(EX248) );
or2  gate( .a(EX242), .b(EX244), .O(EX249) );
or2  gate( .a(EX246), .b(EX249), .O(EX250) );
or2  gate( .a(EX248), .b(EX250), .O(N782) );
nor2 gate300( .a(N754), .b(N755), .O(N785) );
nor2 gate301( .a(N757), .b(N758), .O(N786) );
nor2 gate302( .a(N759), .b(N760), .O(N787) );
inv1 gate( .a(N700),.O(N700_NOT) );
inv1 gate( .a(N773),.O(N773_NOT));
and2 gate( .a(N700_NOT), .b(p101), .O(EX251) );
and2 gate( .a(N773_NOT), .b(EX251), .O(EX252) );
and2 gate( .a(N700), .b(p102), .O(EX253) );
and2 gate( .a(N773_NOT), .b(EX253), .O(EX254) );
and2 gate( .a(N700_NOT), .b(p103), .O(EX255) );
and2 gate( .a(N773), .b(EX255), .O(EX256) );
and2 gate( .a(N700), .b(p104), .O(EX257) );
and2 gate( .a(N773), .b(EX257), .O(EX258) );
or2  gate( .a(EX252), .b(EX254), .O(EX259) );
or2  gate( .a(EX256), .b(EX259), .O(EX260) );
or2  gate( .a(EX258), .b(EX260), .O(N788) );
and2 gate304( .a(N700), .b(N773), .O(N789) );
nor2 gate305( .a(N708), .b(N778), .O(N790) );
and2 gate306( .a(N708), .b(N778), .O(N791) );
nor2 gate307( .a(N717), .b(N782), .O(N792) );
and2 gate308( .a(N717), .b(N782), .O(N793) );
and2 gate309( .a(N219), .b(N786), .O(N794) );
nand2 gate310( .a(N628), .b(N773), .O(N795) );
nand2 gate311( .a(N795), .b(N747), .O(N796) );
nor2 gate312( .a(N788), .b(N789), .O(N802) );
nor2 gate313( .a(N790), .b(N791), .O(N803) );
nor2 gate314( .a(N792), .b(N793), .O(N804) );
nor2 gate315( .a(N340), .b(N794), .O(N805) );
nor2 gate316( .a(N692), .b(N796), .O(N806) );
inv1 gate( .a(N692),.O(N692_NOT) );
inv1 gate( .a(N796),.O(N796_NOT));
and2 gate( .a(N692_NOT), .b(p105), .O(EX261) );
and2 gate( .a(N796_NOT), .b(EX261), .O(EX262) );
and2 gate( .a(N692), .b(p106), .O(EX263) );
and2 gate( .a(N796_NOT), .b(EX263), .O(EX264) );
and2 gate( .a(N692_NOT), .b(p107), .O(EX265) );
and2 gate( .a(N796), .b(EX265), .O(EX266) );
and2 gate( .a(N692), .b(p108), .O(EX267) );
and2 gate( .a(N796), .b(EX267), .O(EX268) );
or2  gate( .a(EX262), .b(EX264), .O(EX269) );
or2  gate( .a(EX266), .b(EX269), .O(EX270) );
or2  gate( .a(EX268), .b(EX270), .O(N807) );
and2 gate318( .a(N219), .b(N802), .O(N808) );
and2 gate319( .a(N219), .b(N803), .O(N809) );
and2 gate320( .a(N219), .b(N804), .O(N810) );
nand4 gate321( .a(N805), .b(N787), .c(N731), .d(N529), .O(N811) );
nand2 gate322( .a(N619), .b(N796), .O(N812) );
nand3 gate323( .a(N609), .b(N619), .c(N796), .O(N813) );
nand4 gate324( .a(N600), .b(N609), .c(N619), .d(N796), .O(N814) );
nand4 gate325( .a(N738), .b(N765), .c(N766), .d(N814), .O(N815) );
nand3 gate326( .a(N741), .b(N764), .c(N813), .O(N819) );
nand2 gate327( .a(N744), .b(N812), .O(N822) );
nor2 gate328( .a(N806), .b(N807), .O(N825) );
inv1 gate( .a(N335),.O(N335_NOT) );
inv1 gate( .a(N808),.O(N808_NOT));
and2 gate( .a(N335_NOT), .b(p109), .O(EX271) );
and2 gate( .a(N808_NOT), .b(EX271), .O(EX272) );
and2 gate( .a(N335), .b(p110), .O(EX273) );
and2 gate( .a(N808_NOT), .b(EX273), .O(EX274) );
and2 gate( .a(N335_NOT), .b(p111), .O(EX275) );
and2 gate( .a(N808), .b(EX275), .O(EX276) );
and2 gate( .a(N335), .b(p112), .O(EX277) );
and2 gate( .a(N808), .b(EX277), .O(EX278) );
or2  gate( .a(EX272), .b(EX274), .O(EX279) );
or2  gate( .a(EX276), .b(EX279), .O(EX280) );
or2  gate( .a(EX278), .b(EX280), .O(N826) );
nor2 gate330( .a(N336), .b(N809), .O(N827) );
nor2 gate331( .a(N338), .b(N810), .O(N828) );
inv1 gate332( .a(N811), .O(N829) );
nor2 gate333( .a(N665), .b(N815), .O(N830) );
and2 gate334( .a(N665), .b(N815), .O(N831) );
nor2 gate335( .a(N673), .b(N819), .O(N832) );
and2 gate336( .a(N673), .b(N819), .O(N833) );
nor2 gate337( .a(N682), .b(N822), .O(N834) );
inv1 gate( .a(N682),.O(N682_NOT) );
inv1 gate( .a(N822),.O(N822_NOT));
and2 gate( .a(N682_NOT), .b(p113), .O(EX281) );
and2 gate( .a(N822_NOT), .b(EX281), .O(EX282) );
and2 gate( .a(N682), .b(p114), .O(EX283) );
and2 gate( .a(N822_NOT), .b(EX283), .O(EX284) );
and2 gate( .a(N682_NOT), .b(p115), .O(EX285) );
and2 gate( .a(N822), .b(EX285), .O(EX286) );
and2 gate( .a(N682), .b(p116), .O(EX287) );
and2 gate( .a(N822), .b(EX287), .O(EX288) );
or2  gate( .a(EX282), .b(EX284), .O(EX289) );
or2  gate( .a(EX286), .b(EX289), .O(EX290) );
or2  gate( .a(EX288), .b(EX290), .O(N835) );
and2 gate339( .a(N219), .b(N825), .O(N836) );
nand3 gate340( .a(N826), .b(N777), .c(N704), .O(N837) );
nand4 gate341( .a(N827), .b(N781), .c(N712), .d(N527), .O(N838) );
nand4 gate342( .a(N828), .b(N785), .c(N721), .d(N528), .O(N839) );
inv1 gate343( .a(N829), .O(N840) );
nand2 gate344( .a(N815), .b(N593), .O(N841) );
nor2 gate345( .a(N830), .b(N831), .O(N842) );
nor2 gate346( .a(N832), .b(N833), .O(N843) );
nor2 gate347( .a(N834), .b(N835), .O(N844) );
nor2 gate348( .a(N334), .b(N836), .O(N845) );
inv1 gate349( .a(N837), .O(N846) );
inv1 gate350( .a(N838), .O(N847) );
inv1 gate351( .a(N839), .O(N848) );
and2 gate352( .a(N735), .b(N841), .O(N849) );
buf1 gate353( .a(N840), .O(N850) );
inv1 gate( .a(N219),.O(N219_NOT) );
inv1 gate( .a(N842),.O(N842_NOT));
and2 gate( .a(N219_NOT), .b(p117), .O(EX291) );
and2 gate( .a(N842_NOT), .b(EX291), .O(EX292) );
and2 gate( .a(N219), .b(p118), .O(EX293) );
and2 gate( .a(N842_NOT), .b(EX293), .O(EX294) );
and2 gate( .a(N219_NOT), .b(p119), .O(EX295) );
and2 gate( .a(N842), .b(EX295), .O(EX296) );
and2 gate( .a(N219), .b(p120), .O(EX297) );
and2 gate( .a(N842), .b(EX297), .O(EX298) );
or2  gate( .a(EX292), .b(EX294), .O(EX299) );
or2  gate( .a(EX296), .b(EX299), .O(EX300) );
or2  gate( .a(EX298), .b(EX300), .O(N851) );
and2 gate355( .a(N219), .b(N843), .O(N852) );
and2 gate356( .a(N219), .b(N844), .O(N853) );
nand3 gate357( .a(N845), .b(N772), .c(N696), .O(N854) );
inv1 gate358( .a(N846), .O(N855) );
inv1 gate359( .a(N847), .O(N856) );
inv1 gate360( .a(N848), .O(N857) );
inv1 gate361( .a(N849), .O(N858) );
inv1 gate( .a(N417),.O(N417_NOT) );
inv1 gate( .a(N851),.O(N851_NOT));
and2 gate( .a(N417_NOT), .b(p121), .O(EX301) );
and2 gate( .a(N851_NOT), .b(EX301), .O(EX302) );
and2 gate( .a(N417), .b(p122), .O(EX303) );
and2 gate( .a(N851_NOT), .b(EX303), .O(EX304) );
and2 gate( .a(N417_NOT), .b(p123), .O(EX305) );
and2 gate( .a(N851), .b(EX305), .O(EX306) );
and2 gate( .a(N417), .b(p124), .O(EX307) );
and2 gate( .a(N851), .b(EX307), .O(EX308) );
or2  gate( .a(EX302), .b(EX304), .O(EX309) );
or2  gate( .a(EX306), .b(EX309), .O(EX310) );
or2  gate( .a(EX308), .b(EX310), .O(N859) );
nor2 gate363( .a(N332), .b(N852), .O(N860) );
nor2 gate364( .a(N333), .b(N853), .O(N861) );
inv1 gate365( .a(N854), .O(N862) );
buf1 gate366( .a(N855), .O(N863) );
buf1 gate367( .a(N856), .O(N864) );
buf1 gate368( .a(N857), .O(N865) );
buf1 gate369( .a(N858), .O(N866) );
nand3 gate370( .a(N859), .b(N769), .c(N669), .O(N867) );
nand3 gate371( .a(N860), .b(N770), .c(N677), .O(N868) );
nand3 gate372( .a(N861), .b(N771), .c(N686), .O(N869) );
inv1 gate373( .a(N862), .O(N870) );
inv1 gate374( .a(N867), .O(N871) );
inv1 gate375( .a(N868), .O(N872) );
inv1 gate376( .a(N869), .O(N873) );
buf1 gate377( .a(N870), .O(N874) );
inv1 gate378( .a(N871), .O(N875) );
inv1 gate379( .a(N872), .O(N876) );
inv1 gate380( .a(N873), .O(N877) );
buf1 gate381( .a(N875), .O(N878) );
buf1 gate382( .a(N876), .O(N879) );
buf1 gate383( .a(N877), .O(N880) );

xor2 gate( .a(X_1), .b(N1_new), .O(N1) );
xor2 gate( .a(X_2), .b(N8_new), .O(N8) );
xor2 gate( .a(X_3), .b(N13_new), .O(N13) );
xor2 gate( .a(X_4), .b(N17_new), .O(N17) );
xor2 gate( .a(X_5), .b(N1_new), .O(N1) );
xor2 gate( .a(X_6), .b(N13_new), .O(N13) );
xor2 gate( .a(X_7), .b(N17_new), .O(N17) );
xor2 gate( .a(X_8), .b(N26_new), .O(N26) );
xor2 gate( .a(X_9), .b(N29_new), .O(N29) );
xor2 gate( .a(X_10), .b(N36_new), .O(N36) );
xor2 gate( .a(X_11), .b(N42_new), .O(N42) );
xor2 gate( .a(X_12), .b(N1_new), .O(N1) );
xor2 gate( .a(X_13), .b(N26_new), .O(N26) );
xor2 gate( .a(X_14), .b(N51_new), .O(N51) );
xor2 gate( .a(X_15), .b(N1_new), .O(N1) );
xor2 gate( .a(X_16), .b(N8_new), .O(N8) );
xor2 gate( .a(X_17), .b(N17_new), .O(N17) );
xor2 gate( .a(X_18), .b(N51_new), .O(N51) );
xor2 gate( .a(X_19), .b(N1_new), .O(N1) );
xor2 gate( .a(X_20), .b(N8_new), .O(N8) );
xor2 gate( .a(X_21), .b(N13_new), .O(N13) );
xor2 gate( .a(X_22), .b(N55_new), .O(N55) );
xor2 gate( .a(X_23), .b(N42_new), .O(N42) );
xor2 gate( .a(X_24), .b(N59_new), .O(N59) );
xor2 gate( .a(X_25), .b(N68_new), .O(N68) );
xor2 gate( .a(X_26), .b(N72_new), .O(N72) );
xor2 gate( .a(X_27), .b(N29_new), .O(N29) );
xor2 gate( .a(X_28), .b(N68_new), .O(N68) );
xor2 gate( .a(X_29), .b(N59_new), .O(N59) );
xor2 gate( .a(X_30), .b(N68_new), .O(N68) );
xor2 gate( .a(X_31), .b(N74_new), .O(N74) );
xor2 gate( .a(X_32), .b(N29_new), .O(N29) );
xor2 gate( .a(X_33), .b(N75_new), .O(N75) );
xor2 gate( .a(X_34), .b(N80_new), .O(N80) );
xor2 gate( .a(X_35), .b(N29_new), .O(N29) );
xor2 gate( .a(X_36), .b(N42_new), .O(N42) );
xor2 gate( .a(X_37), .b(N75_new), .O(N75) );
xor2 gate( .a(X_38), .b(N29_new), .O(N29) );
xor2 gate( .a(X_39), .b(N36_new), .O(N36) );
xor2 gate( .a(X_40), .b(N80_new), .O(N80) );
xor2 gate( .a(X_41), .b(N29_new), .O(N29) );
xor2 gate( .a(X_42), .b(N36_new), .O(N36) );
xor2 gate( .a(X_43), .b(N42_new), .O(N42) );
xor2 gate( .a(X_44), .b(N59_new), .O(N59) );
xor2 gate( .a(X_45), .b(N75_new), .O(N75) );
xor2 gate( .a(X_46), .b(N80_new), .O(N80) );
xor2 gate( .a(X_47), .b(N42_new), .O(N42) );
xor2 gate( .a(X_48), .b(N59_new), .O(N59) );
xor2 gate( .a(X_49), .b(N75_new), .O(N75) );
xor2 gate( .a(X_50), .b(N36_new), .O(N36) );
xor2 gate( .a(X_51), .b(N59_new), .O(N59) );
xor2 gate( .a(X_52), .b(N80_new), .O(N80) );
xor2 gate( .a(X_53), .b(N36_new), .O(N36) );
xor2 gate( .a(X_54), .b(N42_new), .O(N42) );
xor2 gate( .a(X_55), .b(N59_new), .O(N59) );
xor2 gate( .a(X_56), .b(N85_new), .O(N85) );
xor2 gate( .a(X_57), .b(N86_new), .O(N86) );
xor2 gate( .a(X_58), .b(N87_new), .O(N87) );
xor2 gate( .a(X_59), .b(N88_new), .O(N88) );
xor2 gate( .a(X_60), .b(N91_new), .O(N91) );
xor2 gate( .a(X_61), .b(N96_new), .O(N96) );
xor2 gate( .a(X_62), .b(N91_new), .O(N91) );
xor2 gate( .a(X_63), .b(N96_new), .O(N96) );
xor2 gate( .a(X_64), .b(N101_new), .O(N101) );
xor2 gate( .a(X_65), .b(N106_new), .O(N106) );
xor2 gate( .a(X_66), .b(N101_new), .O(N101) );
xor2 gate( .a(X_67), .b(N106_new), .O(N106) );
xor2 gate( .a(X_68), .b(N101_new), .O(N101) );
xor2 gate( .a(X_69), .b(N106_new), .O(N106) );
xor2 gate( .a(X_70), .b(N101_new), .O(N101) );
xor2 gate( .a(X_71), .b(N106_new), .O(N106) );
xor2 gate( .a(X_72), .b(N111_new), .O(N111) );
xor2 gate( .a(X_73), .b(N116_new), .O(N116) );
xor2 gate( .a(X_74), .b(N111_new), .O(N111) );
xor2 gate( .a(X_75), .b(N116_new), .O(N116) );
xor2 gate( .a(X_76), .b(N111_new), .O(N111) );
xor2 gate( .a(X_77), .b(N116_new), .O(N116) );
xor2 gate( .a(X_78), .b(N111_new), .O(N111) );
xor2 gate( .a(X_79), .b(N116_new), .O(N116) );
xor2 gate( .a(X_80), .b(N121_new), .O(N121) );
xor2 gate( .a(X_81), .b(N126_new), .O(N126) );
xor2 gate( .a(X_82), .b(N121_new), .O(N121) );
xor2 gate( .a(X_83), .b(N126_new), .O(N126) );
xor2 gate( .a(X_84), .b(N8_new), .O(N8) );
xor2 gate( .a(X_85), .b(N138_new), .O(N138) );
xor2 gate( .a(X_86), .b(N268_new), .O(N268) );
xor2 gate( .a(X_87), .b(N51_new), .O(N51) );
xor2 gate( .a(X_88), .b(N138_new), .O(N138) );
xor2 gate( .a(X_89), .b(N17_new), .O(N17) );
xor2 gate( .a(X_90), .b(N138_new), .O(N138) );
xor2 gate( .a(X_91), .b(N138_new), .O(N138) );
xor2 gate( .a(X_92), .b(N152_new), .O(N152) );
xor2 gate( .a(X_93), .b(N59_new), .O(N59) );
xor2 gate( .a(X_94), .b(N156_new), .O(N156) );
xor2 gate( .a(X_95), .b(N17_new), .O(N17) );
xor2 gate( .a(X_96), .b(N42_new), .O(N42) );
xor2 gate( .a(X_97), .b(N17_new), .O(N17) );
xor2 gate( .a(X_98), .b(N42_new), .O(N42) );
xor2 gate( .a(X_99), .b(N159_new), .O(N159) );
xor2 gate( .a(X_100), .b(N165_new), .O(N165) );
xor2 gate( .a(X_101), .b(N159_new), .O(N159) );
xor2 gate( .a(X_102), .b(N165_new), .O(N165) );
xor2 gate( .a(X_103), .b(N159_new), .O(N159) );
xor2 gate( .a(X_104), .b(N165_new), .O(N165) );
xor2 gate( .a(X_105), .b(N159_new), .O(N159) );
xor2 gate( .a(X_106), .b(N165_new), .O(N165) );
xor2 gate( .a(X_107), .b(N171_new), .O(N171) );
xor2 gate( .a(X_108), .b(N177_new), .O(N177) );
xor2 gate( .a(X_109), .b(N171_new), .O(N171) );
xor2 gate( .a(X_110), .b(N177_new), .O(N177) );
xor2 gate( .a(X_111), .b(N171_new), .O(N171) );
xor2 gate( .a(X_112), .b(N177_new), .O(N177) );
xor2 gate( .a(X_113), .b(N171_new), .O(N171) );
xor2 gate( .a(X_114), .b(N177_new), .O(N177) );
xor2 gate( .a(X_115), .b(N183_new), .O(N183) );
xor2 gate( .a(X_116), .b(N189_new), .O(N189) );
xor2 gate( .a(X_117), .b(N183_new), .O(N183) );
xor2 gate( .a(X_118), .b(N189_new), .O(N189) );
xor2 gate( .a(X_119), .b(N195_new), .O(N195) );
xor2 gate( .a(X_120), .b(N201_new), .O(N201) );
xor2 gate( .a(X_121), .b(N195_new), .O(N195) );
xor2 gate( .a(X_122), .b(N201_new), .O(N201) );
xor2 gate( .a(X_123), .b(N91_new), .O(N91) );
xor2 gate( .a(X_124), .b(N210_new), .O(N210) );
xor2 gate( .a(X_125), .b(N96_new), .O(N96) );
xor2 gate( .a(X_126), .b(N210_new), .O(N210) );
xor2 gate( .a(X_127), .b(N101_new), .O(N101) );
xor2 gate( .a(X_128), .b(N210_new), .O(N210) );
xor2 gate( .a(X_129), .b(N106_new), .O(N106) );
xor2 gate( .a(X_130), .b(N210_new), .O(N210) );
xor2 gate( .a(X_131), .b(N111_new), .O(N111) );
xor2 gate( .a(X_132), .b(N210_new), .O(N210) );
xor2 gate( .a(X_133), .b(N255_new), .O(N255) );
xor2 gate( .a(X_134), .b(N259_new), .O(N259) );
xor2 gate( .a(X_135), .b(N255_new), .O(N255) );
xor2 gate( .a(X_136), .b(N259_new), .O(N259) );
xor2 gate( .a(X_137), .b(N255_new), .O(N255) );
xor2 gate( .a(X_138), .b(N259_new), .O(N259) );
xor2 gate( .a(X_139), .b(N116_new), .O(N116) );
xor2 gate( .a(X_140), .b(N210_new), .O(N210) );
xor2 gate( .a(X_141), .b(N255_new), .O(N255) );
xor2 gate( .a(X_142), .b(N260_new), .O(N260) );
xor2 gate( .a(X_143), .b(N121_new), .O(N121) );
xor2 gate( .a(X_144), .b(N210_new), .O(N210) );
xor2 gate( .a(X_145), .b(N255_new), .O(N255) );
xor2 gate( .a(X_146), .b(N267_new), .O(N267) );
xor2 gate( .a(X_147), .b(N89_new), .O(N89) );
xor2 gate( .a(X_148), .b(N90_new), .O(N90) );
xor2 gate( .a(X_149), .b(N388), .O(N388_new) );
xor2 gate( .a(X_150), .b(N389), .O(N389_new) );
xor2 gate( .a(X_151), .b(N390), .O(N390_new) );
xor2 gate( .a(X_152), .b(N391), .O(N391_new) );
xor2 gate( .a(X_153), .b(N73_new), .O(N73) );
xor2 gate( .a(X_154), .b(N210_new), .O(N210) );
xor2 gate( .a(X_155), .b(N418), .O(N418_new) );
xor2 gate( .a(X_156), .b(N419), .O(N419_new) );
xor2 gate( .a(X_157), .b(N420), .O(N420_new) );
xor2 gate( .a(X_158), .b(N421), .O(N421_new) );
xor2 gate( .a(X_159), .b(N422), .O(N422_new) );
xor2 gate( .a(X_160), .b(N423), .O(N423_new) );
xor2 gate( .a(X_161), .b(N55_new), .O(N55) );
xor2 gate( .a(X_162), .b(N17_new), .O(N17) );
xor2 gate( .a(X_163), .b(N55_new), .O(N55) );
xor2 gate( .a(X_164), .b(N59_new), .O(N59) );
xor2 gate( .a(X_165), .b(N156_new), .O(N156) );
xor2 gate( .a(X_166), .b(N17_new), .O(N17) );
xor2 gate( .a(X_167), .b(N446), .O(N446_new) );
xor2 gate( .a(X_168), .b(N447), .O(N447_new) );
xor2 gate( .a(X_169), .b(N448), .O(N448_new) );
xor2 gate( .a(X_170), .b(N449), .O(N449_new) );
xor2 gate( .a(X_171), .b(N450), .O(N450_new) );
xor2 gate( .a(X_172), .b(N143_new), .O(N143) );
xor2 gate( .a(X_173), .b(N146_new), .O(N146) );
xor2 gate( .a(X_174), .b(N149_new), .O(N149) );
xor2 gate( .a(X_175), .b(N153_new), .O(N153) );
xor2 gate( .a(X_176), .b(N1_new), .O(N1) );
xor2 gate( .a(X_177), .b(N130_new), .O(N130) );
xor2 gate( .a(X_178), .b(N130_new), .O(N130) );
xor2 gate( .a(X_179), .b(N130_new), .O(N130) );
xor2 gate( .a(X_180), .b(N130_new), .O(N130) );
xor2 gate( .a(X_181), .b(N130_new), .O(N130) );
xor2 gate( .a(X_182), .b(N130_new), .O(N130) );
xor2 gate( .a(X_183), .b(N135_new), .O(N135) );
xor2 gate( .a(X_184), .b(N135_new), .O(N135) );
xor2 gate( .a(X_185), .b(N135_new), .O(N135) );
xor2 gate( .a(X_186), .b(N135_new), .O(N135) );
xor2 gate( .a(X_187), .b(N91_new), .O(N91) );
xor2 gate( .a(X_188), .b(N91_new), .O(N91) );
xor2 gate( .a(X_189), .b(N91_new), .O(N91) );
xor2 gate( .a(X_190), .b(N96_new), .O(N96) );
xor2 gate( .a(X_191), .b(N96_new), .O(N96) );
xor2 gate( .a(X_192), .b(N96_new), .O(N96) );
xor2 gate( .a(X_193), .b(N101_new), .O(N101) );
xor2 gate( .a(X_194), .b(N106_new), .O(N106) );
xor2 gate( .a(X_195), .b(N143_new), .O(N143) );
xor2 gate( .a(X_196), .b(N111_new), .O(N111) );
xor2 gate( .a(X_197), .b(N146_new), .O(N146) );
xor2 gate( .a(X_198), .b(N116_new), .O(N116) );
xor2 gate( .a(X_199), .b(N149_new), .O(N149) );
xor2 gate( .a(X_200), .b(N121_new), .O(N121) );
xor2 gate( .a(X_201), .b(N153_new), .O(N153) );
xor2 gate( .a(X_202), .b(N126_new), .O(N126) );
xor2 gate( .a(X_203), .b(N130_new), .O(N130) );
xor2 gate( .a(X_204), .b(N130_new), .O(N130) );
xor2 gate( .a(X_205), .b(N207_new), .O(N207) );
xor2 gate( .a(X_206), .b(N207_new), .O(N207) );
xor2 gate( .a(X_207), .b(N159_new), .O(N159) );
xor2 gate( .a(X_208), .b(N165_new), .O(N165) );
xor2 gate( .a(X_209), .b(N171_new), .O(N171) );
xor2 gate( .a(X_210), .b(N171_new), .O(N171) );
xor2 gate( .a(X_211), .b(N171_new), .O(N171) );
xor2 gate( .a(X_212), .b(N177_new), .O(N177) );
xor2 gate( .a(X_213), .b(N183_new), .O(N183) );
xor2 gate( .a(X_214), .b(N189_new), .O(N189) );
xor2 gate( .a(X_215), .b(N195_new), .O(N195) );
xor2 gate( .a(X_216), .b(N201_new), .O(N201) );
xor2 gate( .a(X_217), .b(N159_new), .O(N159) );
xor2 gate( .a(X_218), .b(N159_new), .O(N159) );
xor2 gate( .a(X_219), .b(N246_new), .O(N246) );
xor2 gate( .a(X_220), .b(N165_new), .O(N165) );
xor2 gate( .a(X_221), .b(N165_new), .O(N165) );
xor2 gate( .a(X_222), .b(N246_new), .O(N246) );
xor2 gate( .a(X_223), .b(N246_new), .O(N246) );
xor2 gate( .a(X_224), .b(N246_new), .O(N246) );
xor2 gate( .a(X_225), .b(N171_new), .O(N171) );
xor2 gate( .a(X_226), .b(N171_new), .O(N171) );
xor2 gate( .a(X_227), .b(N246_new), .O(N246) );
xor2 gate( .a(X_228), .b(N177_new), .O(N177) );
xor2 gate( .a(X_229), .b(N177_new), .O(N177) );
xor2 gate( .a(X_230), .b(N246_new), .O(N246) );
xor2 gate( .a(X_231), .b(N183_new), .O(N183) );
xor2 gate( .a(X_232), .b(N183_new), .O(N183) );
xor2 gate( .a(X_233), .b(N246_new), .O(N246) );
xor2 gate( .a(X_234), .b(N246_new), .O(N246) );
xor2 gate( .a(X_235), .b(N246_new), .O(N246) );
xor2 gate( .a(X_236), .b(N189_new), .O(N189) );
xor2 gate( .a(X_237), .b(N189_new), .O(N189) );
xor2 gate( .a(X_238), .b(N246_new), .O(N246) );
xor2 gate( .a(X_239), .b(N195_new), .O(N195) );
xor2 gate( .a(X_240), .b(N195_new), .O(N195) );
xor2 gate( .a(X_241), .b(N246_new), .O(N246) );
xor2 gate( .a(X_242), .b(N201_new), .O(N201) );
xor2 gate( .a(X_243), .b(N201_new), .O(N201) );
xor2 gate( .a(X_244), .b(N246_new), .O(N246) );
xor2 gate( .a(X_245), .b(N261_new), .O(N261) );
xor2 gate( .a(X_246), .b(N261_new), .O(N261) );
xor2 gate( .a(X_247), .b(N261_new), .O(N261) );
xor2 gate( .a(X_248), .b(N228_new), .O(N228) );
xor2 gate( .a(X_249), .b(N237_new), .O(N237) );
xor2 gate( .a(X_250), .b(N228_new), .O(N228) );
xor2 gate( .a(X_251), .b(N237_new), .O(N237) );
xor2 gate( .a(X_252), .b(N228_new), .O(N228) );
xor2 gate( .a(X_253), .b(N237_new), .O(N237) );
xor2 gate( .a(X_254), .b(N228_new), .O(N228) );
xor2 gate( .a(X_255), .b(N237_new), .O(N237) );
xor2 gate( .a(X_256), .b(N228_new), .O(N228) );
xor2 gate( .a(X_257), .b(N237_new), .O(N237) );
xor2 gate( .a(X_258), .b(N228_new), .O(N228) );
xor2 gate( .a(X_259), .b(N228_new), .O(N228) );
xor2 gate( .a(X_260), .b(N228_new), .O(N228) );
xor2 gate( .a(X_261), .b(N237_new), .O(N237) );
xor2 gate( .a(X_262), .b(N228_new), .O(N228) );
xor2 gate( .a(X_263), .b(N237_new), .O(N237) );
xor2 gate( .a(X_264), .b(N261_new), .O(N261) );
xor2 gate( .a(X_265), .b(N261_new), .O(N261) );
xor2 gate( .a(X_266), .b(N228_new), .O(N228) );
xor2 gate( .a(X_267), .b(N237_new), .O(N237) );
xor2 gate( .a(X_268), .b(N767), .O(N767_new) );
xor2 gate( .a(X_269), .b(N768), .O(N768_new) );
xor2 gate( .a(X_270), .b(N219_new), .O(N219) );
xor2 gate( .a(X_271), .b(N219_new), .O(N219) );
xor2 gate( .a(X_272), .b(N219_new), .O(N219) );
xor2 gate( .a(X_273), .b(N219_new), .O(N219) );
xor2 gate( .a(X_274), .b(N219_new), .O(N219) );
xor2 gate( .a(X_275), .b(N850), .O(N850_new) );
xor2 gate( .a(X_276), .b(N219_new), .O(N219) );
xor2 gate( .a(X_277), .b(N219_new), .O(N219) );
xor2 gate( .a(X_278), .b(N219_new), .O(N219) );
xor2 gate( .a(X_279), .b(N219_new), .O(N219) );
xor2 gate( .a(X_280), .b(N219_new), .O(N219) );
xor2 gate( .a(X_281), .b(N863), .O(N863_new) );
xor2 gate( .a(X_282), .b(N864), .O(N864_new) );
xor2 gate( .a(X_283), .b(N865), .O(N865_new) );
xor2 gate( .a(X_284), .b(N866), .O(N866_new) );
xor2 gate( .a(X_285), .b(N874), .O(N874_new) );
xor2 gate( .a(X_286), .b(N878), .O(N878_new) );
xor2 gate( .a(X_287), .b(N879), .O(N879_new) );
xor2 gate( .a(X_288), .b(N880), .O(N880_new) );
endmodule