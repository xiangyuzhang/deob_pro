
module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);

input N1_new,N5_new,N9_new,N13_new,N17_new,N21_new,N25_new,N29_new,N33_new,N37_new,
      N41_new,N45_new,N49_new,N53_new,N57_new,N61_new,N65_new,N69_new,N73_new,N77_new,
      N81_new,N85_new,N89_new,N93_new,N97_new,N101_new,N105_new,N109_new,N113_new,N117_new,
      N121_new,N125_new,N129_new,N130_new,N131_new,N132_new,N133_new,N134_new,N135_new,N136_new,
      N137_new;

input p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,
        p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,
        p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,
        p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,
        p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,
        p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,
        p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,
        p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,
        p81,p82,p83,p84,X_1,X_2,X_3,X_4,X_5,X_6,X_7,X_8,X_9,X_10,X_11,X_12,X_13,X_14,X_15,X_16,X_17,X_18,X_19,X_20,X_21,X_22,X_23,X_24,X_25,X_26,X_27,X_28,X_29,X_30,X_31,X_32,X_33,X_34,X_35,X_36,X_37,X_38,X_39,X_40,X_41,X_42,X_43,X_44,X_45,X_46,X_47,X_48,X_49,X_50,X_51,X_52,X_53,X_54,X_55,X_56,X_57,X_58,X_59,X_60,X_61,X_62,X_63,X_64,X_65,X_66,X_67,X_68,X_69,X_70,X_71,X_72,X_73,X_74,X_75,X_76,X_77,X_78,X_79,X_80,X_81,X_82,X_83,X_84,X_85,X_86,X_87,X_88,X_89,X_90,X_91,X_92,X_93,X_94,X_95,X_96,X_97,X_98,X_99,X_100,X_101,X_102,X_103,X_104,X_105,X_106,X_107,X_108,X_109,X_110,X_111,X_112,X_113,X_114,X_115,X_116,X_117,X_118,X_119,X_120,X_121,X_122,X_123,X_124,X_125,X_126,X_127,X_128,X_129,X_130,X_131,X_132,X_133,X_134,X_135,X_136,X_137,X_138,X_139,X_140,X_141,X_142,X_143,X_144,X_145,X_146,X_147,X_148,X_149,X_150,X_151,X_152,X_153,X_154,X_155,X_156,X_157,X_158,X_159,X_160,X_161,X_162,X_163,X_164,X_165,X_166,X_167,X_168,X_169,X_170,X_171,X_172,X_173,X_174,X_175,X_176,X_177,X_178;

output N724_new,N725_new,N726_new,N727_new,N728_new,N729_new,N730_new,N731_new,N732_new,N733_new,
       N734_new,N735_new,N736_new,N737_new,N738_new,N739_new,N740_new,N741_new,N742_new,N743_new,
       N744_new,N745_new,N746_new,N747_new,N748_new,N749_new,N750_new,N751_new,N752_new,N753_new,
       N754_new,N755_new;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,
     N65_NOT,N69_NOT,N73_NOT,N77_NOT,N81_NOT,N85_NOT,N97_NOT,N101_NOT,N131_NOT,N137_NOT,
     N135_NOT,N137_NOT,N256_NOT,N257_NOT,N278_NOT,N279_NOT,N282_NOT,N283_NOT,N288_NOT,N289_NOT,
     N302_NOT,N305_NOT,N272_NOT,N340_NOT,N321_NOT,N353_NOT,N419_NOT,N650_NOT,N445_NOT,N650_NOT,
     N419_NOT,N655_NOT,N5_NOT,N693_NOT,N13_NOT,N695_NOT,N41_NOT,N702_NOT,N77_NOT,N711_NOT,
     N97_NOT,N716_NOT,EX1,EX2,EX3,EX4,EX5,EX6,EX7,EX8,EX9,EX10,
     EX11,EX12,EX13,EX14,EX15,EX16,EX17,EX18,EX19,EX20,
     EX21,EX22,EX23,EX24,EX25,EX26,EX27,EX28,EX29,EX30,
     EX31,EX32,EX33,EX34,EX35,EX36,EX37,EX38,EX39,EX40,
     EX41,EX42,EX43,EX44,EX45,EX46,EX47,EX48,EX49,EX50,
     EX51,EX52,EX53,EX54,EX55,EX56,EX57,EX58,EX59,EX60,
     EX61,EX62,EX63,EX64,EX65,EX66,EX67,EX68,EX69,EX70,
     EX71,EX72,EX73,EX74,EX75,EX76,EX77,EX78,EX79,EX80,
     EX81,EX82,EX83,EX84,EX85,EX86,EX87,EX88,EX89,EX90,
     EX91,EX92,EX93,EX94,EX95,EX96,EX97,EX98,EX99,EX100,
     EX101,EX102,EX103,EX104,EX105,EX106,EX107,EX108,EX109,EX110,
     EX111,EX112,EX113,EX114,EX115,EX116,EX117,EX118,EX119,EX120,
     EX121,EX122,EX123,EX124,EX125,EX126,EX127,EX128,EX129,EX130,
     EX131,EX132,EX133,EX134,EX135,EX136,EX137,EX138,EX139,EX140,
     EX141,EX142,EX143,EX144,EX145,EX146,EX147,EX148,EX149,EX150,
     EX151,EX152,EX153,EX154,EX155,EX156,EX157,EX158,EX159,EX160,
     EX161,EX162,EX163,EX164,EX165,EX166,EX167,EX168,EX169,EX170,
     EX171,EX172,EX173,EX174,EX175,EX176,EX177,EX178,EX179,EX180,
     EX181,EX182,EX183,EX184,EX185,EX186,EX187,EX188,EX189,EX190,
     EX191,EX192,EX193,EX194,EX195,EX196,EX197,EX198,EX199,EX200,
     EX201,EX202,EX203,EX204,EX205,EX206,EX207,EX208,EX209,EX210,N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755;


xor2 gate1( .a(N1), .b(N5), .O(N250) );
xor2 gate2( .a(N9), .b(N13), .O(N251) );
xor2 gate3( .a(N17), .b(N21), .O(N252) );
xor2 gate4( .a(N25), .b(N29), .O(N253) );
xor2 gate5( .a(N33), .b(N37), .O(N254) );
xor2 gate6( .a(N41), .b(N45), .O(N255) );
xor2 gate7( .a(N49), .b(N53), .O(N256) );
xor2 gate8( .a(N57), .b(N61), .O(N257) );
inv1 gate( .a(N65),.O(N65_NOT) );
inv1 gate( .a(N69),.O(N69_NOT));
and2 gate( .a(N65_NOT), .b(p1), .O(EX1) );
and2 gate( .a(N69_NOT), .b(EX1), .O(EX2) );
and2 gate( .a(N65), .b(p2), .O(EX3) );
and2 gate( .a(N69_NOT), .b(EX3), .O(EX4) );
and2 gate( .a(N65_NOT), .b(p3), .O(EX5) );
and2 gate( .a(N69), .b(EX5), .O(EX6) );
and2 gate( .a(N65), .b(p4), .O(EX7) );
and2 gate( .a(N69), .b(EX7), .O(EX8) );
or2  gate( .a(EX2), .b(EX4), .O(EX9) );
or2  gate( .a(EX6), .b(EX9), .O(EX10) );
or2  gate( .a(EX8), .b(EX10), .O(N258) );
inv1 gate( .a(N73),.O(N73_NOT) );
inv1 gate( .a(N77),.O(N77_NOT));
and2 gate( .a(N73_NOT), .b(p5), .O(EX11) );
and2 gate( .a(N77_NOT), .b(EX11), .O(EX12) );
and2 gate( .a(N73), .b(p6), .O(EX13) );
and2 gate( .a(N77_NOT), .b(EX13), .O(EX14) );
and2 gate( .a(N73_NOT), .b(p7), .O(EX15) );
and2 gate( .a(N77), .b(EX15), .O(EX16) );
and2 gate( .a(N73), .b(p8), .O(EX17) );
and2 gate( .a(N77), .b(EX17), .O(EX18) );
or2  gate( .a(EX12), .b(EX14), .O(EX19) );
or2  gate( .a(EX16), .b(EX19), .O(EX20) );
or2  gate( .a(EX18), .b(EX20), .O(N259) );
inv1 gate( .a(N81),.O(N81_NOT) );
inv1 gate( .a(N85),.O(N85_NOT));
and2 gate( .a(N81_NOT), .b(p9), .O(EX21) );
and2 gate( .a(N85_NOT), .b(EX21), .O(EX22) );
and2 gate( .a(N81), .b(p10), .O(EX23) );
and2 gate( .a(N85_NOT), .b(EX23), .O(EX24) );
and2 gate( .a(N81_NOT), .b(p11), .O(EX25) );
and2 gate( .a(N85), .b(EX25), .O(EX26) );
and2 gate( .a(N81), .b(p12), .O(EX27) );
and2 gate( .a(N85), .b(EX27), .O(EX28) );
or2  gate( .a(EX22), .b(EX24), .O(EX29) );
or2  gate( .a(EX26), .b(EX29), .O(EX30) );
or2  gate( .a(EX28), .b(EX30), .O(N260) );
xor2 gate12( .a(N89), .b(N93), .O(N261) );
inv1 gate( .a(N97),.O(N97_NOT) );
inv1 gate( .a(N101),.O(N101_NOT));
and2 gate( .a(N97_NOT), .b(p13), .O(EX31) );
and2 gate( .a(N101_NOT), .b(EX31), .O(EX32) );
and2 gate( .a(N97), .b(p14), .O(EX33) );
and2 gate( .a(N101_NOT), .b(EX33), .O(EX34) );
and2 gate( .a(N97_NOT), .b(p15), .O(EX35) );
and2 gate( .a(N101), .b(EX35), .O(EX36) );
and2 gate( .a(N97), .b(p16), .O(EX37) );
and2 gate( .a(N101), .b(EX37), .O(EX38) );
or2  gate( .a(EX32), .b(EX34), .O(EX39) );
or2  gate( .a(EX36), .b(EX39), .O(EX40) );
or2  gate( .a(EX38), .b(EX40), .O(N262) );
xor2 gate14( .a(N105), .b(N109), .O(N263) );
xor2 gate15( .a(N113), .b(N117), .O(N264) );
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
inv1 gate( .a(N131),.O(N131_NOT) );
inv1 gate( .a(N137),.O(N137_NOT));
and2 gate( .a(N131_NOT), .b(p17), .O(EX41) );
and2 gate( .a(N137_NOT), .b(EX41), .O(EX42) );
and2 gate( .a(N131), .b(p18), .O(EX43) );
and2 gate( .a(N137_NOT), .b(EX43), .O(EX44) );
and2 gate( .a(N131_NOT), .b(p19), .O(EX45) );
and2 gate( .a(N137), .b(EX45), .O(EX46) );
and2 gate( .a(N131), .b(p20), .O(EX47) );
and2 gate( .a(N137), .b(EX47), .O(EX48) );
or2  gate( .a(EX42), .b(EX44), .O(EX49) );
or2  gate( .a(EX46), .b(EX49), .O(EX50) );
or2  gate( .a(EX48), .b(EX50), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
inv1 gate( .a(N135),.O(N135_NOT) );
inv1 gate( .a(N137),.O(N137_NOT));
and2 gate( .a(N135_NOT), .b(p21), .O(EX51) );
and2 gate( .a(N137_NOT), .b(EX51), .O(EX52) );
and2 gate( .a(N135), .b(p22), .O(EX53) );
and2 gate( .a(N137_NOT), .b(EX53), .O(EX54) );
and2 gate( .a(N135_NOT), .b(p23), .O(EX55) );
and2 gate( .a(N137), .b(EX55), .O(EX56) );
and2 gate( .a(N135), .b(p24), .O(EX57) );
and2 gate( .a(N137), .b(EX57), .O(EX58) );
or2  gate( .a(EX52), .b(EX54), .O(EX59) );
or2  gate( .a(EX56), .b(EX59), .O(EX60) );
or2  gate( .a(EX58), .b(EX60), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );
xor2 gate26( .a(N33), .b(N49), .O(N275) );
xor2 gate27( .a(N5), .b(N21), .O(N276) );
xor2 gate28( .a(N37), .b(N53), .O(N277) );
xor2 gate29( .a(N9), .b(N25), .O(N278) );
xor2 gate30( .a(N41), .b(N57), .O(N279) );
xor2 gate31( .a(N13), .b(N29), .O(N280) );
xor2 gate32( .a(N45), .b(N61), .O(N281) );
xor2 gate33( .a(N65), .b(N81), .O(N282) );
xor2 gate34( .a(N97), .b(N113), .O(N283) );
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );
xor2 gate37( .a(N73), .b(N89), .O(N286) );
xor2 gate38( .a(N105), .b(N121), .O(N287) );
xor2 gate39( .a(N77), .b(N93), .O(N288) );
xor2 gate40( .a(N109), .b(N125), .O(N289) );
xor2 gate41( .a(N250), .b(N251), .O(N290) );
xor2 gate42( .a(N252), .b(N253), .O(N293) );
xor2 gate43( .a(N254), .b(N255), .O(N296) );
inv1 gate( .a(N256),.O(N256_NOT) );
inv1 gate( .a(N257),.O(N257_NOT));
and2 gate( .a(N256_NOT), .b(p25), .O(EX61) );
and2 gate( .a(N257_NOT), .b(EX61), .O(EX62) );
and2 gate( .a(N256), .b(p26), .O(EX63) );
and2 gate( .a(N257_NOT), .b(EX63), .O(EX64) );
and2 gate( .a(N256_NOT), .b(p27), .O(EX65) );
and2 gate( .a(N257), .b(EX65), .O(EX66) );
and2 gate( .a(N256), .b(p28), .O(EX67) );
and2 gate( .a(N257), .b(EX67), .O(EX68) );
or2  gate( .a(EX62), .b(EX64), .O(EX69) );
or2  gate( .a(EX66), .b(EX69), .O(EX70) );
or2  gate( .a(EX68), .b(EX70), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );
xor2 gate46( .a(N260), .b(N261), .O(N305) );
xor2 gate47( .a(N262), .b(N263), .O(N308) );
xor2 gate48( .a(N264), .b(N265), .O(N311) );
xor2 gate49( .a(N274), .b(N275), .O(N314) );
xor2 gate50( .a(N276), .b(N277), .O(N315) );
inv1 gate( .a(N278),.O(N278_NOT) );
inv1 gate( .a(N279),.O(N279_NOT));
and2 gate( .a(N278_NOT), .b(p29), .O(EX71) );
and2 gate( .a(N279_NOT), .b(EX71), .O(EX72) );
and2 gate( .a(N278), .b(p30), .O(EX73) );
and2 gate( .a(N279_NOT), .b(EX73), .O(EX74) );
and2 gate( .a(N278_NOT), .b(p31), .O(EX75) );
and2 gate( .a(N279), .b(EX75), .O(EX76) );
and2 gate( .a(N278), .b(p32), .O(EX77) );
and2 gate( .a(N279), .b(EX77), .O(EX78) );
or2  gate( .a(EX72), .b(EX74), .O(EX79) );
or2  gate( .a(EX76), .b(EX79), .O(EX80) );
or2  gate( .a(EX78), .b(EX80), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );
inv1 gate( .a(N282),.O(N282_NOT) );
inv1 gate( .a(N283),.O(N283_NOT));
and2 gate( .a(N282_NOT), .b(p33), .O(EX81) );
and2 gate( .a(N283_NOT), .b(EX81), .O(EX82) );
and2 gate( .a(N282), .b(p34), .O(EX83) );
and2 gate( .a(N283_NOT), .b(EX83), .O(EX84) );
and2 gate( .a(N282_NOT), .b(p35), .O(EX85) );
and2 gate( .a(N283), .b(EX85), .O(EX86) );
and2 gate( .a(N282), .b(p36), .O(EX87) );
and2 gate( .a(N283), .b(EX87), .O(EX88) );
or2  gate( .a(EX82), .b(EX84), .O(EX89) );
or2  gate( .a(EX86), .b(EX89), .O(EX90) );
or2  gate( .a(EX88), .b(EX90), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );
xor2 gate55( .a(N286), .b(N287), .O(N320) );
inv1 gate( .a(N288),.O(N288_NOT) );
inv1 gate( .a(N289),.O(N289_NOT));
and2 gate( .a(N288_NOT), .b(p37), .O(EX91) );
and2 gate( .a(N289_NOT), .b(EX91), .O(EX92) );
and2 gate( .a(N288), .b(p38), .O(EX93) );
and2 gate( .a(N289_NOT), .b(EX93), .O(EX94) );
and2 gate( .a(N288_NOT), .b(p39), .O(EX95) );
and2 gate( .a(N289), .b(EX95), .O(EX96) );
and2 gate( .a(N288), .b(p40), .O(EX97) );
and2 gate( .a(N289), .b(EX97), .O(EX98) );
or2  gate( .a(EX92), .b(EX94), .O(EX99) );
or2  gate( .a(EX96), .b(EX99), .O(EX100) );
or2  gate( .a(EX98), .b(EX100), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );
xor2 gate58( .a(N296), .b(N299), .O(N339) );
xor2 gate59( .a(N290), .b(N296), .O(N340) );
xor2 gate60( .a(N293), .b(N299), .O(N341) );
inv1 gate( .a(N302),.O(N302_NOT) );
inv1 gate( .a(N305),.O(N305_NOT));
and2 gate( .a(N302_NOT), .b(p41), .O(EX101) );
and2 gate( .a(N305_NOT), .b(EX101), .O(EX102) );
and2 gate( .a(N302), .b(p42), .O(EX103) );
and2 gate( .a(N305_NOT), .b(EX103), .O(EX104) );
and2 gate( .a(N302_NOT), .b(p43), .O(EX105) );
and2 gate( .a(N305), .b(EX105), .O(EX106) );
and2 gate( .a(N302), .b(p44), .O(EX107) );
and2 gate( .a(N305), .b(EX107), .O(EX108) );
or2  gate( .a(EX102), .b(EX104), .O(EX109) );
or2  gate( .a(EX106), .b(EX109), .O(EX110) );
or2  gate( .a(EX108), .b(EX110), .O(N342) );
xor2 gate62( .a(N308), .b(N311), .O(N343) );
xor2 gate63( .a(N302), .b(N308), .O(N344) );
xor2 gate64( .a(N305), .b(N311), .O(N345) );
xor2 gate65( .a(N266), .b(N342), .O(N346) );
xor2 gate66( .a(N267), .b(N343), .O(N347) );
xor2 gate67( .a(N268), .b(N344), .O(N348) );
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );
xor2 gate70( .a(N271), .b(N339), .O(N351) );
inv1 gate( .a(N272),.O(N272_NOT) );
inv1 gate( .a(N340),.O(N340_NOT));
and2 gate( .a(N272_NOT), .b(p45), .O(EX111) );
and2 gate( .a(N340_NOT), .b(EX111), .O(EX112) );
and2 gate( .a(N272), .b(p46), .O(EX113) );
and2 gate( .a(N340_NOT), .b(EX113), .O(EX114) );
and2 gate( .a(N272_NOT), .b(p47), .O(EX115) );
and2 gate( .a(N340), .b(EX115), .O(EX116) );
and2 gate( .a(N272), .b(p48), .O(EX117) );
and2 gate( .a(N340), .b(EX117), .O(EX118) );
or2  gate( .a(EX112), .b(EX114), .O(EX119) );
or2  gate( .a(EX116), .b(EX119), .O(EX120) );
or2  gate( .a(EX118), .b(EX120), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );
xor2 gate74( .a(N315), .b(N347), .O(N367) );
xor2 gate75( .a(N316), .b(N348), .O(N380) );
xor2 gate76( .a(N317), .b(N349), .O(N393) );
xor2 gate77( .a(N318), .b(N350), .O(N406) );
xor2 gate78( .a(N319), .b(N351), .O(N419) );
xor2 gate79( .a(N320), .b(N352), .O(N432) );
inv1 gate( .a(N321),.O(N321_NOT) );
inv1 gate( .a(N353),.O(N353_NOT));
and2 gate( .a(N321_NOT), .b(p49), .O(EX121) );
and2 gate( .a(N353_NOT), .b(EX121), .O(EX122) );
and2 gate( .a(N321), .b(p50), .O(EX123) );
and2 gate( .a(N353_NOT), .b(EX123), .O(EX124) );
and2 gate( .a(N321_NOT), .b(p51), .O(EX125) );
and2 gate( .a(N353), .b(EX125), .O(EX126) );
and2 gate( .a(N321), .b(p52), .O(EX127) );
and2 gate( .a(N353), .b(EX127), .O(EX128) );
or2  gate( .a(EX122), .b(EX124), .O(EX129) );
or2  gate( .a(EX126), .b(EX129), .O(EX130) );
or2  gate( .a(EX128), .b(EX130), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
inv1 gate( .a(N419),.O(N419_NOT) );
inv1 gate( .a(N650),.O(N650_NOT));
and2 gate( .a(N419_NOT), .b(p53), .O(EX131) );
and2 gate( .a(N650_NOT), .b(EX131), .O(EX132) );
and2 gate( .a(N419), .b(p54), .O(EX133) );
and2 gate( .a(N650_NOT), .b(EX133), .O(EX134) );
and2 gate( .a(N419_NOT), .b(p55), .O(EX135) );
and2 gate( .a(N650), .b(EX135), .O(EX136) );
and2 gate( .a(N419), .b(p56), .O(EX137) );
and2 gate( .a(N650), .b(EX137), .O(EX138) );
or2  gate( .a(EX132), .b(EX134), .O(EX139) );
or2  gate( .a(EX136), .b(EX139), .O(EX140) );
or2  gate( .a(EX138), .b(EX140), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
inv1 gate( .a(N445),.O(N445_NOT) );
inv1 gate( .a(N650),.O(N650_NOT));
and2 gate( .a(N445_NOT), .b(p57), .O(EX141) );
and2 gate( .a(N650_NOT), .b(EX141), .O(EX142) );
and2 gate( .a(N445), .b(p58), .O(EX143) );
and2 gate( .a(N650_NOT), .b(EX143), .O(EX144) );
and2 gate( .a(N445_NOT), .b(p59), .O(EX145) );
and2 gate( .a(N650), .b(EX145), .O(EX146) );
and2 gate( .a(N445), .b(p60), .O(EX147) );
and2 gate( .a(N650), .b(EX147), .O(EX148) );
or2  gate( .a(EX142), .b(EX144), .O(EX149) );
or2  gate( .a(EX146), .b(EX149), .O(EX150) );
or2  gate( .a(EX148), .b(EX150), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
inv1 gate( .a(N419),.O(N419_NOT) );
inv1 gate( .a(N655),.O(N655_NOT));
and2 gate( .a(N419_NOT), .b(p61), .O(EX151) );
and2 gate( .a(N655_NOT), .b(EX151), .O(EX152) );
and2 gate( .a(N419), .b(p62), .O(EX153) );
and2 gate( .a(N655_NOT), .b(EX153), .O(EX154) );
and2 gate( .a(N419_NOT), .b(p63), .O(EX155) );
and2 gate( .a(N655), .b(EX155), .O(EX156) );
and2 gate( .a(N419), .b(p64), .O(EX157) );
and2 gate( .a(N655), .b(EX157), .O(EX158) );
or2  gate( .a(EX152), .b(EX154), .O(EX159) );
or2  gate( .a(EX156), .b(EX159), .O(EX160) );
or2  gate( .a(EX158), .b(EX160), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );
inv1 gate( .a(N5),.O(N5_NOT) );
inv1 gate( .a(N693),.O(N693_NOT));
and2 gate( .a(N5_NOT), .b(p65), .O(EX161) );
and2 gate( .a(N693_NOT), .b(EX161), .O(EX162) );
and2 gate( .a(N5), .b(p66), .O(EX163) );
and2 gate( .a(N693_NOT), .b(EX163), .O(EX164) );
and2 gate( .a(N5_NOT), .b(p67), .O(EX165) );
and2 gate( .a(N693), .b(EX165), .O(EX166) );
and2 gate( .a(N5), .b(p68), .O(EX167) );
and2 gate( .a(N693), .b(EX167), .O(EX168) );
or2  gate( .a(EX162), .b(EX164), .O(EX169) );
or2  gate( .a(EX166), .b(EX169), .O(EX170) );
or2  gate( .a(EX168), .b(EX170), .O(N725) );
xor2 gate173( .a(N9), .b(N694), .O(N726) );
inv1 gate( .a(N13),.O(N13_NOT) );
inv1 gate( .a(N695),.O(N695_NOT));
and2 gate( .a(N13_NOT), .b(p69), .O(EX171) );
and2 gate( .a(N695_NOT), .b(EX171), .O(EX172) );
and2 gate( .a(N13), .b(p70), .O(EX173) );
and2 gate( .a(N695_NOT), .b(EX173), .O(EX174) );
and2 gate( .a(N13_NOT), .b(p71), .O(EX175) );
and2 gate( .a(N695), .b(EX175), .O(EX176) );
and2 gate( .a(N13), .b(p72), .O(EX177) );
and2 gate( .a(N695), .b(EX177), .O(EX178) );
or2  gate( .a(EX172), .b(EX174), .O(EX179) );
or2  gate( .a(EX176), .b(EX179), .O(EX180) );
or2  gate( .a(EX178), .b(EX180), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );
xor2 gate176( .a(N21), .b(N697), .O(N729) );
xor2 gate177( .a(N25), .b(N698), .O(N730) );
xor2 gate178( .a(N29), .b(N699), .O(N731) );
xor2 gate179( .a(N33), .b(N700), .O(N732) );
xor2 gate180( .a(N37), .b(N701), .O(N733) );
inv1 gate( .a(N41),.O(N41_NOT) );
inv1 gate( .a(N702),.O(N702_NOT));
and2 gate( .a(N41_NOT), .b(p73), .O(EX181) );
and2 gate( .a(N702_NOT), .b(EX181), .O(EX182) );
and2 gate( .a(N41), .b(p74), .O(EX183) );
and2 gate( .a(N702_NOT), .b(EX183), .O(EX184) );
and2 gate( .a(N41_NOT), .b(p75), .O(EX185) );
and2 gate( .a(N702), .b(EX185), .O(EX186) );
and2 gate( .a(N41), .b(p76), .O(EX187) );
and2 gate( .a(N702), .b(EX187), .O(EX188) );
or2  gate( .a(EX182), .b(EX184), .O(EX189) );
or2  gate( .a(EX186), .b(EX189), .O(EX190) );
or2  gate( .a(EX188), .b(EX190), .O(N734) );
xor2 gate182( .a(N45), .b(N703), .O(N735) );
xor2 gate183( .a(N49), .b(N704), .O(N736) );
xor2 gate184( .a(N53), .b(N705), .O(N737) );
xor2 gate185( .a(N57), .b(N706), .O(N738) );
xor2 gate186( .a(N61), .b(N707), .O(N739) );
xor2 gate187( .a(N65), .b(N708), .O(N740) );
xor2 gate188( .a(N69), .b(N709), .O(N741) );
xor2 gate189( .a(N73), .b(N710), .O(N742) );
inv1 gate( .a(N77),.O(N77_NOT) );
inv1 gate( .a(N711),.O(N711_NOT));
and2 gate( .a(N77_NOT), .b(p77), .O(EX191) );
and2 gate( .a(N711_NOT), .b(EX191), .O(EX192) );
and2 gate( .a(N77), .b(p78), .O(EX193) );
and2 gate( .a(N711_NOT), .b(EX193), .O(EX194) );
and2 gate( .a(N77_NOT), .b(p79), .O(EX195) );
and2 gate( .a(N711), .b(EX195), .O(EX196) );
and2 gate( .a(N77), .b(p80), .O(EX197) );
and2 gate( .a(N711), .b(EX197), .O(EX198) );
or2  gate( .a(EX192), .b(EX194), .O(EX199) );
or2  gate( .a(EX196), .b(EX199), .O(EX200) );
or2  gate( .a(EX198), .b(EX200), .O(N743) );
xor2 gate191( .a(N81), .b(N712), .O(N744) );
xor2 gate192( .a(N85), .b(N713), .O(N745) );
xor2 gate193( .a(N89), .b(N714), .O(N746) );
xor2 gate194( .a(N93), .b(N715), .O(N747) );
inv1 gate( .a(N97),.O(N97_NOT) );
inv1 gate( .a(N716),.O(N716_NOT));
and2 gate( .a(N97_NOT), .b(p81), .O(EX201) );
and2 gate( .a(N716_NOT), .b(EX201), .O(EX202) );
and2 gate( .a(N97), .b(p82), .O(EX203) );
and2 gate( .a(N716_NOT), .b(EX203), .O(EX204) );
and2 gate( .a(N97_NOT), .b(p83), .O(EX205) );
and2 gate( .a(N716), .b(EX205), .O(EX206) );
and2 gate( .a(N97), .b(p84), .O(EX207) );
and2 gate( .a(N716), .b(EX207), .O(EX208) );
or2  gate( .a(EX202), .b(EX204), .O(EX209) );
or2  gate( .a(EX206), .b(EX209), .O(EX210) );
or2  gate( .a(EX208), .b(EX210), .O(N748) );
xor2 gate196( .a(N101), .b(N717), .O(N749) );
xor2 gate197( .a(N105), .b(N718), .O(N750) );
xor2 gate198( .a(N109), .b(N719), .O(N751) );
xor2 gate199( .a(N113), .b(N720), .O(N752) );
xor2 gate200( .a(N117), .b(N721), .O(N753) );
xor2 gate201( .a(N121), .b(N722), .O(N754) );
xor2 gate202( .a(N125), .b(N723), .O(N755) );

xor2 gate( .a(X_1), .b(N1_new), .O(N1) );
xor2 gate( .a(X_2), .b(N5_new), .O(N5) );
xor2 gate( .a(X_3), .b(N9_new), .O(N9) );
xor2 gate( .a(X_4), .b(N13_new), .O(N13) );
xor2 gate( .a(X_5), .b(N17_new), .O(N17) );
xor2 gate( .a(X_6), .b(N21_new), .O(N21) );
xor2 gate( .a(X_7), .b(N25_new), .O(N25) );
xor2 gate( .a(X_8), .b(N29_new), .O(N29) );
xor2 gate( .a(X_9), .b(N33_new), .O(N33) );
xor2 gate( .a(X_10), .b(N37_new), .O(N37) );
xor2 gate( .a(X_11), .b(N41_new), .O(N41) );
xor2 gate( .a(X_12), .b(N45_new), .O(N45) );
xor2 gate( .a(X_13), .b(N49_new), .O(N49) );
xor2 gate( .a(X_14), .b(N53_new), .O(N53) );
xor2 gate( .a(X_15), .b(N57_new), .O(N57) );
xor2 gate( .a(X_16), .b(N61_new), .O(N61) );
xor2 gate( .a(X_17), .b(N65_new), .O(N65) );
xor2 gate( .a(X_18), .b(N69_new), .O(N69) );
xor2 gate( .a(X_19), .b(N65_new), .O(N65) );
xor2 gate( .a(X_20), .b(N69_new), .O(N69) );
xor2 gate( .a(X_21), .b(N65_new), .O(N65) );
xor2 gate( .a(X_22), .b(N69_new), .O(N69) );
xor2 gate( .a(X_23), .b(N73_new), .O(N73) );
xor2 gate( .a(X_24), .b(N77_new), .O(N77) );
xor2 gate( .a(X_25), .b(N73_new), .O(N73) );
xor2 gate( .a(X_26), .b(N77_new), .O(N77) );
xor2 gate( .a(X_27), .b(N73_new), .O(N73) );
xor2 gate( .a(X_28), .b(N77_new), .O(N77) );
xor2 gate( .a(X_29), .b(N81_new), .O(N81) );
xor2 gate( .a(X_30), .b(N85_new), .O(N85) );
xor2 gate( .a(X_31), .b(N81_new), .O(N81) );
xor2 gate( .a(X_32), .b(N85_new), .O(N85) );
xor2 gate( .a(X_33), .b(N81_new), .O(N81) );
xor2 gate( .a(X_34), .b(N85_new), .O(N85) );
xor2 gate( .a(X_35), .b(N89_new), .O(N89) );
xor2 gate( .a(X_36), .b(N93_new), .O(N93) );
xor2 gate( .a(X_37), .b(N97_new), .O(N97) );
xor2 gate( .a(X_38), .b(N101_new), .O(N101) );
xor2 gate( .a(X_39), .b(N97_new), .O(N97) );
xor2 gate( .a(X_40), .b(N101_new), .O(N101) );
xor2 gate( .a(X_41), .b(N97_new), .O(N97) );
xor2 gate( .a(X_42), .b(N101_new), .O(N101) );
xor2 gate( .a(X_43), .b(N105_new), .O(N105) );
xor2 gate( .a(X_44), .b(N109_new), .O(N109) );
xor2 gate( .a(X_45), .b(N113_new), .O(N113) );
xor2 gate( .a(X_46), .b(N117_new), .O(N117) );
xor2 gate( .a(X_47), .b(N121_new), .O(N121) );
xor2 gate( .a(X_48), .b(N125_new), .O(N125) );
xor2 gate( .a(X_49), .b(N129_new), .O(N129) );
xor2 gate( .a(X_50), .b(N137_new), .O(N137) );
xor2 gate( .a(X_51), .b(N130_new), .O(N130) );
xor2 gate( .a(X_52), .b(N137_new), .O(N137) );
xor2 gate( .a(X_53), .b(N131_new), .O(N131) );
xor2 gate( .a(X_54), .b(N137_new), .O(N137) );
xor2 gate( .a(X_55), .b(N131_new), .O(N131) );
xor2 gate( .a(X_56), .b(N137_new), .O(N137) );
xor2 gate( .a(X_57), .b(N131_new), .O(N131) );
xor2 gate( .a(X_58), .b(N137_new), .O(N137) );
xor2 gate( .a(X_59), .b(N132_new), .O(N132) );
xor2 gate( .a(X_60), .b(N137_new), .O(N137) );
xor2 gate( .a(X_61), .b(N133_new), .O(N133) );
xor2 gate( .a(X_62), .b(N137_new), .O(N137) );
xor2 gate( .a(X_63), .b(N134_new), .O(N134) );
xor2 gate( .a(X_64), .b(N137_new), .O(N137) );
xor2 gate( .a(X_65), .b(N135_new), .O(N135) );
xor2 gate( .a(X_66), .b(N137_new), .O(N137) );
xor2 gate( .a(X_67), .b(N135_new), .O(N135) );
xor2 gate( .a(X_68), .b(N137_new), .O(N137) );
xor2 gate( .a(X_69), .b(N135_new), .O(N135) );
xor2 gate( .a(X_70), .b(N137_new), .O(N137) );
xor2 gate( .a(X_71), .b(N136_new), .O(N136) );
xor2 gate( .a(X_72), .b(N137_new), .O(N137) );
xor2 gate( .a(X_73), .b(N1_new), .O(N1) );
xor2 gate( .a(X_74), .b(N17_new), .O(N17) );
xor2 gate( .a(X_75), .b(N33_new), .O(N33) );
xor2 gate( .a(X_76), .b(N49_new), .O(N49) );
xor2 gate( .a(X_77), .b(N5_new), .O(N5) );
xor2 gate( .a(X_78), .b(N21_new), .O(N21) );
xor2 gate( .a(X_79), .b(N37_new), .O(N37) );
xor2 gate( .a(X_80), .b(N53_new), .O(N53) );
xor2 gate( .a(X_81), .b(N9_new), .O(N9) );
xor2 gate( .a(X_82), .b(N25_new), .O(N25) );
xor2 gate( .a(X_83), .b(N41_new), .O(N41) );
xor2 gate( .a(X_84), .b(N57_new), .O(N57) );
xor2 gate( .a(X_85), .b(N13_new), .O(N13) );
xor2 gate( .a(X_86), .b(N29_new), .O(N29) );
xor2 gate( .a(X_87), .b(N45_new), .O(N45) );
xor2 gate( .a(X_88), .b(N61_new), .O(N61) );
xor2 gate( .a(X_89), .b(N65_new), .O(N65) );
xor2 gate( .a(X_90), .b(N81_new), .O(N81) );
xor2 gate( .a(X_91), .b(N97_new), .O(N97) );
xor2 gate( .a(X_92), .b(N113_new), .O(N113) );
xor2 gate( .a(X_93), .b(N69_new), .O(N69) );
xor2 gate( .a(X_94), .b(N85_new), .O(N85) );
xor2 gate( .a(X_95), .b(N101_new), .O(N101) );
xor2 gate( .a(X_96), .b(N117_new), .O(N117) );
xor2 gate( .a(X_97), .b(N73_new), .O(N73) );
xor2 gate( .a(X_98), .b(N89_new), .O(N89) );
xor2 gate( .a(X_99), .b(N105_new), .O(N105) );
xor2 gate( .a(X_100), .b(N121_new), .O(N121) );
xor2 gate( .a(X_101), .b(N77_new), .O(N77) );
xor2 gate( .a(X_102), .b(N93_new), .O(N93) );
xor2 gate( .a(X_103), .b(N109_new), .O(N109) );
xor2 gate( .a(X_104), .b(N125_new), .O(N125) );
xor2 gate( .a(X_105), .b(N724), .O(N724_new) );
xor2 gate( .a(X_106), .b(N1_new), .O(N1) );
xor2 gate( .a(X_107), .b(N5_new), .O(N5) );
xor2 gate( .a(X_108), .b(N5_new), .O(N5) );
xor2 gate( .a(X_109), .b(N5_new), .O(N5) );
xor2 gate( .a(X_110), .b(N725), .O(N725_new) );
xor2 gate( .a(X_111), .b(N726), .O(N726_new) );
xor2 gate( .a(X_112), .b(N9_new), .O(N9) );
xor2 gate( .a(X_113), .b(N13_new), .O(N13) );
xor2 gate( .a(X_114), .b(N13_new), .O(N13) );
xor2 gate( .a(X_115), .b(N13_new), .O(N13) );
xor2 gate( .a(X_116), .b(N727), .O(N727_new) );
xor2 gate( .a(X_117), .b(N728), .O(N728_new) );
xor2 gate( .a(X_118), .b(N17_new), .O(N17) );
xor2 gate( .a(X_119), .b(N729), .O(N729_new) );
xor2 gate( .a(X_120), .b(N21_new), .O(N21) );
xor2 gate( .a(X_121), .b(N730), .O(N730_new) );
xor2 gate( .a(X_122), .b(N25_new), .O(N25) );
xor2 gate( .a(X_123), .b(N731), .O(N731_new) );
xor2 gate( .a(X_124), .b(N29_new), .O(N29) );
xor2 gate( .a(X_125), .b(N732), .O(N732_new) );
xor2 gate( .a(X_126), .b(N33_new), .O(N33) );
xor2 gate( .a(X_127), .b(N733), .O(N733_new) );
xor2 gate( .a(X_128), .b(N37_new), .O(N37) );
xor2 gate( .a(X_129), .b(N41_new), .O(N41) );
xor2 gate( .a(X_130), .b(N41_new), .O(N41) );
xor2 gate( .a(X_131), .b(N41_new), .O(N41) );
xor2 gate( .a(X_132), .b(N734), .O(N734_new) );
xor2 gate( .a(X_133), .b(N735), .O(N735_new) );
xor2 gate( .a(X_134), .b(N45_new), .O(N45) );
xor2 gate( .a(X_135), .b(N736), .O(N736_new) );
xor2 gate( .a(X_136), .b(N49_new), .O(N49) );
xor2 gate( .a(X_137), .b(N737), .O(N737_new) );
xor2 gate( .a(X_138), .b(N53_new), .O(N53) );
xor2 gate( .a(X_139), .b(N738), .O(N738_new) );
xor2 gate( .a(X_140), .b(N57_new), .O(N57) );
xor2 gate( .a(X_141), .b(N739), .O(N739_new) );
xor2 gate( .a(X_142), .b(N61_new), .O(N61) );
xor2 gate( .a(X_143), .b(N740), .O(N740_new) );
xor2 gate( .a(X_144), .b(N65_new), .O(N65) );
xor2 gate( .a(X_145), .b(N741), .O(N741_new) );
xor2 gate( .a(X_146), .b(N69_new), .O(N69) );
xor2 gate( .a(X_147), .b(N742), .O(N742_new) );
xor2 gate( .a(X_148), .b(N73_new), .O(N73) );
xor2 gate( .a(X_149), .b(N77_new), .O(N77) );
xor2 gate( .a(X_150), .b(N77_new), .O(N77) );
xor2 gate( .a(X_151), .b(N77_new), .O(N77) );
xor2 gate( .a(X_152), .b(N743), .O(N743_new) );
xor2 gate( .a(X_153), .b(N744), .O(N744_new) );
xor2 gate( .a(X_154), .b(N81_new), .O(N81) );
xor2 gate( .a(X_155), .b(N745), .O(N745_new) );
xor2 gate( .a(X_156), .b(N85_new), .O(N85) );
xor2 gate( .a(X_157), .b(N746), .O(N746_new) );
xor2 gate( .a(X_158), .b(N89_new), .O(N89) );
xor2 gate( .a(X_159), .b(N747), .O(N747_new) );
xor2 gate( .a(X_160), .b(N93_new), .O(N93) );
xor2 gate( .a(X_161), .b(N97_new), .O(N97) );
xor2 gate( .a(X_162), .b(N97_new), .O(N97) );
xor2 gate( .a(X_163), .b(N97_new), .O(N97) );
xor2 gate( .a(X_164), .b(N748), .O(N748_new) );
xor2 gate( .a(X_165), .b(N749), .O(N749_new) );
xor2 gate( .a(X_166), .b(N101_new), .O(N101) );
xor2 gate( .a(X_167), .b(N750), .O(N750_new) );
xor2 gate( .a(X_168), .b(N105_new), .O(N105) );
xor2 gate( .a(X_169), .b(N751), .O(N751_new) );
xor2 gate( .a(X_170), .b(N109_new), .O(N109) );
xor2 gate( .a(X_171), .b(N752), .O(N752_new) );
xor2 gate( .a(X_172), .b(N113_new), .O(N113) );
xor2 gate( .a(X_173), .b(N753), .O(N753_new) );
xor2 gate( .a(X_174), .b(N117_new), .O(N117) );
xor2 gate( .a(X_175), .b(N754), .O(N754_new) );
xor2 gate( .a(X_176), .b(N121_new), .O(N121) );
xor2 gate( .a(X_177), .b(N755), .O(N755_new) );
xor2 gate( .a(X_178), .b(N125_new), .O(N125) );
endmodule