module	c17 (N1,N2,N3,N4,N5,N6,N7,N8,N9,N12,N13,N14);
input N1,N2,N3,N4,N5 //RE__PI;

input D_0,D_1,D_2,D_3,D_4,D_5,D_6,D_7 //RE__ALLOW(00,01,10,11);
output N6,N7;
wire N9,N12,N13,N14,D_0_NOT,D_1_NOT,MUX_O_0,ED_0,ED_1,ED_2,ED_3,ED_4,ED_5,ED_6,ED_7,ED_8,ED_9,D_2_NOT,D_3_NOT,MUX_O_1,ED_10,ED_11,ED_12,ED_13,ED_14,ED_15,ED_16,ED_17,ED_18,ED_19,D_4_NOT,D_5_NOT,MUX_O_2,ED_20,ED_21,ED_22,ED_23,ED_24,ED_25,ED_26,ED_27,ED_28,ED_29,D_6_NOT,D_7_NOT,MUX_O_3,ED_30,ED_31,ED_32,ED_33,ED_34,ED_35,ED_36,ED_37,ED_38,ED_39;
nand2 gate1( .a(N1), .b(N3), .O(N14) );
nand2 gate2( .a(N3), .b(N4), .O(N9) );
nand2 gate3( .a(N2), .b(MUX_O_1), .O(N13) );
nand2 gate4( .a(N5), .b(MUX_O_1), .O(N12) );
nand2 gate5( .a(MUX_O_0), .b(MUX_O_3), .O(N6) );
nand2 gate6( .a(N12), .b(N12), .O(N7) );
inv1 gate( .a(D_0),.O(D_0_NOT) );
inv1 gate( .a(D_1),.O(D_1_NOT) );
and2 gate( .a(N1), .b(D_0_NOT), .O(ED_0) );
and2 gate( .a(N14), .b(D_0), .O(ED_1) );
and2 gate( .a(N4), .b(D_0_NOT), .O(ED_2) );
and2 gate( .a(N14), .b(D_0), .O(ED_3) );
and2 gate( .a(ED_0), .b(D_1_NOT), .O(ED_4) );
and2 gate( .a(ED_1), .b(D_1), .O(ED_5) );
and2 gate( .a(ED_2), .b(D_1_NOT), .O(ED_6) );
and2 gate( .a(ED_3), .b(D_1), .O(ED_7) );
or2  gate( .a(ED_4), .b(ED_5), .O(ED_8) );
or2  gate( .a(ED_6), .b(ED_8), .O(ED_9) );
or2  gate( .a(ED_9), .b(ED_7), .O(MUX_O_0) );
inv1 gate( .a(D_2),.O(D_2_NOT) );
inv1 gate( .a(D_3),.O(D_3_NOT) );
and2 gate( .a(N1), .b(D_2_NOT), .O(ED_10) );
and2 gate( .a(N9), .b(D_2), .O(ED_11) );
and2 gate( .a(N4), .b(D_2_NOT), .O(ED_12) );
and2 gate( .a(N9), .b(D_2), .O(ED_13) );
and2 gate( .a(ED_10), .b(D_3_NOT), .O(ED_14) );
and2 gate( .a(ED_11), .b(D_3), .O(ED_15) );
and2 gate( .a(ED_12), .b(D_3_NOT), .O(ED_16) );
and2 gate( .a(ED_13), .b(D_3), .O(ED_17) );
or2  gate( .a(ED_14), .b(ED_15), .O(ED_18) );
or2  gate( .a(ED_16), .b(ED_18), .O(ED_19) );
or2  gate( .a(ED_19), .b(ED_17), .O(MUX_O_1) );
inv1 gate( .a(D_4),.O(D_4_NOT) );
inv1 gate( .a(D_5),.O(D_5_NOT) );
and2 gate( .a(N1), .b(D_4_NOT), .O(ED_20) );
and2 gate( .a(N9), .b(D_4), .O(ED_21) );
and2 gate( .a(N4), .b(D_4_NOT), .O(ED_22) );
and2 gate( .a(N9), .b(D_4), .O(ED_23) );
and2 gate( .a(ED_20), .b(D_5_NOT), .O(ED_24) );
and2 gate( .a(ED_21), .b(D_5), .O(ED_25) );
and2 gate( .a(ED_22), .b(D_5_NOT), .O(ED_26) );
and2 gate( .a(ED_23), .b(D_5), .O(ED_27) );
or2  gate( .a(ED_24), .b(ED_25), .O(ED_28) );
or2  gate( .a(ED_26), .b(ED_28), .O(ED_29) );
or2  gate( .a(ED_29), .b(ED_27), .O(MUX_O_2) );
inv1 gate( .a(D_6),.O(D_6_NOT) );
inv1 gate( .a(D_7),.O(D_7_NOT) );
and2 gate( .a(N1), .b(D_6_NOT), .O(ED_30) );
and2 gate( .a(N13), .b(D_6), .O(ED_31) );
and2 gate( .a(N4), .b(D_6_NOT), .O(ED_32) );
and2 gate( .a(N13), .b(D_6), .O(ED_33) );
and2 gate( .a(ED_30), .b(D_7_NOT), .O(ED_34) );
and2 gate( .a(ED_31), .b(D_7), .O(ED_35) );
and2 gate( .a(ED_32), .b(D_7_NOT), .O(ED_36) );
and2 gate( .a(ED_33), .b(D_7), .O(ED_37) );
or2  gate( .a(ED_34), .b(ED_35), .O(ED_38) );
or2  gate( .a(ED_36), .b(ED_38), .O(ED_39) );
or2  gate( .a(ED_39), .b(ED_37), .O(MUX_O_3) );
endmodule