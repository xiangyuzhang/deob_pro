
module c880 (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
             N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
             N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
             N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
             N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
             N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
             N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
             N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
             N865,N866,N874,N878,N879,N880);

input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;

input p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,
        p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,
        p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,
        p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,
        p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,
        p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,
        p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,
        p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,
        p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,
        p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,
        p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,
        p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,
        p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,
        p131,p132,p133,p134,p135,p136,p137,p138,p139,p140,
        p141,p142,p143,p144,p145,p146,p147,p148,p149,p150,
        p151,p152,p153,p154,p155,p156,p157,p158,p159,p160,
        p161,p162,p163,p164,p165,p166,p167,p168,p169,p170,
        p171,p172,p173,p174,p175,p176,p177,p178,p179,p180,
        p181,p182,p183,p184,p185,p186,p187,p188,p189,p190,
        p191,p192,p193,p194,p195,p196,p197,p198,p199,p200,
        p201,p202,p203,p204,p205,p206,p207,p208,p209,p210,
        p211,p212,p213,p214,p215,p216,p217,p218,p219,p220,
        p221,p222,p223,p224,p225,p226,p227,p228,p229,p230,
        p231,p232,p233,p234,p235,p236,p237,p238,p239,p240,
        p241,p242,p243,p244,p245,p246,p247,p248,p249,p250,
        p251,p252,p253,p254,p255,p256,p257,p258,p259,p260,
        p261,p262,p263,p264,p265,p266,p267,p268,p269,p270,
        p271,p272,p273,p274,p275,p276,p277,p278,p279,p280,
        p281,p282,p283,p284,p285,p286,p287,p288,p289,p290,
        p291,p292,p293,p294,p295,p296,p297,p298,p299,p300,
        p301,p302,p303,p304,p305,p306,p307,p308,p309,p310,
        p311,p312,p313,p314,p315,p316,p317,p318,p319,p320,
        p321,p322,p323,p324,p325,p326,p327,p328,p329,p330,
        p331,p332,p333,p334,p335,p336,p337,p338,p339,p340,
        p341,p342,p343,p344,p345,p346,p347,p348,p349,p350,
        p351,p352,p353,p354,p355,p356,p357,p358,p359,p360,
        p361,p362,p363,p364,p365,p366,p367,p368,p369,p370,
        p371,p372,p373,p374,p375,p376,p377,p378,p379,p380,
        p381,p382,p383,p384,p385,p386,p387,p388,p389,p390,
        p391,p392,p393,p394,p395,p396,p397,p398,p399,p400,
        p401,p402,p403,p404,p405,p406,p407,p408,p409,p410,
        p411,p412,p413,p414,p415,p416,p417,p418,p419,p420,
        p421,p422,p423,p424,p425,p426,p427,p428,p429,p430,
        p431,p432,p433,p434,p435,p436,p437,p438,p439,p440,
        p441,p442,p443,p444;

output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880;

wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,
     N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,
     N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,
     N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,
     N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
     N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
     N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,
     N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
     N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
     N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,
     N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,
     N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,
     N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,
     N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
     N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
     N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
     N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,
     N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,
     N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,
     N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,
     N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,
     N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,
     N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,
     N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
     N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
     N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
     N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
     N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,
     N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,
     N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,
     N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,
     N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
     N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
     N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,
     N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,
     N870,N871,N872,N873,N875,N876,N877,
     N101_NOT,N106_NOT,N101_NOT,N106_NOT,N111_NOT,N116_NOT,N121_NOT,N126_NOT,N17_NOT,N138_NOT,
     N152_NOT,N138_NOT,N17_NOT,N42_NOT,N159_NOT,N165_NOT,N171_NOT,N177_NOT,N171_NOT,N177_NOT,
     N210_NOT,N96_NOT,N210_NOT,N111_NOT,N255_NOT,N259_NOT,N210_NOT,N116_NOT,N255_NOT,N267_NOT,
     N270_NOT,N273_NOT,N280_NOT,N286_NOT,N305_NOT,N306_NOT,N307_NOT,N308_NOT,N322_NOT,N323_NOT,
     N326_NOT,N327_NOT,N330_NOT,N331_NOT,N348_NOT,N73_NOT,N357_NOT,N360_NOT,N363_NOT,N366_NOT,
     N210_NOT,N369_NOT,N407_NOT,N408_NOT,N411_NOT,N412_NOT,N442_NOT,N410_NOT,N143_NOT,N427_NOT,
     N310_NOT,N432_NOT,N443_NOT,N1_NOT,N369_NOT,N437_NOT,N130_NOT,N460_NOT,N130_NOT,N460_NOT,
     N463_NOT,N135_NOT,N91_NOT,N466_NOT,N475_NOT,N476_NOT,N96_NOT,N466_NOT,N477_NOT,N478_NOT,
     N101_NOT,N466_NOT,N146_NOT,N483_NOT,N116_NOT,N466_NOT,N153_NOT,N483_NOT,N130_NOT,N492_NOT,
     N495_NOT,N207_NOT,N451_NOT,N165_NOT,N451_NOT,N171_NOT,N451_NOT,N177_NOT,N451_NOT,N195_NOT,
     N498_NOT,N499_NOT,N317_NOT,N506_NOT,N510_NOT,N511_NOT,N514_NOT,N515_NOT,N516_NOT,N517_NOT,
     N518_NOT,N519_NOT,N488_NOT,N540_NOT,N550_NOT,N551_NOT,N585_NOT,N586_NOT,N553_NOT,N159_NOT,
     N553_NOT,N159_NOT,N557_NOT,N165_NOT,N246_NOT,N557_NOT,N561_NOT,N171_NOT,N565_NOT,N177_NOT,
     N569_NOT,N183_NOT,N569_NOT,N183_NOT,N246_NOT,N569_NOT,N573_NOT,N189_NOT,N581_NOT,N201_NOT,
     N246_NOT,N581_NOT,N587_NOT,N589_NOT,N593_NOT,N590_NOT,N596_NOT,N522_NOT,N609_NOT,N606_NOT,
     N631_NOT,N526_NOT,N635_NOT,N632_NOT,N654_NOT,N651_NOT,N228_NOT,N665_NOT,N237_NOT,N662_NOT,
     N228_NOT,N682_NOT,N237_NOT,N678_NOT,N237_NOT,N687_NOT,N228_NOT,N700_NOT,N228_NOT,N708_NOT,
     N237_NOT,N713_NOT,N228_NOT,N727_NOT,N600_NOT,N678_NOT,N736_NOT,N737_NOT,N748_NOT,N749_NOT,
     N751_NOT,N752_NOT,N756_NOT,N732_NOT,N754_NOT,N755_NOT,N700_NOT,N773_NOT,N700_NOT,N773_NOT,
     N708_NOT,N778_NOT,N628_NOT,N773_NOT,N795_NOT,N747_NOT,N788_NOT,N789_NOT,N792_NOT,N793_NOT,
     N340_NOT,N794_NOT,N692_NOT,N796_NOT,N692_NOT,N796_NOT,N335_NOT,N808_NOT,N665_NOT,N815_NOT,
     N665_NOT,N815_NOT,N682_NOT,N822_NOT,N815_NOT,N593_NOT,N832_NOT,N833_NOT,N219_NOT,N842_NOT,
     N417_NOT,N851_NOT,EX1,EX2,EX3,EX4,EX5,EX6,EX7,EX8,EX9,EX10,
     EX11,EX12,EX13,EX14,EX15,EX16,EX17,EX18,EX19,EX20,
     EX21,EX22,EX23,EX24,EX25,EX26,EX27,EX28,EX29,EX30,
     EX31,EX32,EX33,EX34,EX35,EX36,EX37,EX38,EX39,EX40,
     EX41,EX42,EX43,EX44,EX45,EX46,EX47,EX48,EX49,EX50,
     EX51,EX52,EX53,EX54,EX55,EX56,EX57,EX58,EX59,EX60,
     EX61,EX62,EX63,EX64,EX65,EX66,EX67,EX68,EX69,EX70,
     EX71,EX72,EX73,EX74,EX75,EX76,EX77,EX78,EX79,EX80,
     EX81,EX82,EX83,EX84,EX85,EX86,EX87,EX88,EX89,EX90,
     EX91,EX92,EX93,EX94,EX95,EX96,EX97,EX98,EX99,EX100,
     EX101,EX102,EX103,EX104,EX105,EX106,EX107,EX108,EX109,EX110,
     EX111,EX112,EX113,EX114,EX115,EX116,EX117,EX118,EX119,EX120,
     EX121,EX122,EX123,EX124,EX125,EX126,EX127,EX128,EX129,EX130,
     EX131,EX132,EX133,EX134,EX135,EX136,EX137,EX138,EX139,EX140,
     EX141,EX142,EX143,EX144,EX145,EX146,EX147,EX148,EX149,EX150,
     EX151,EX152,EX153,EX154,EX155,EX156,EX157,EX158,EX159,EX160,
     EX161,EX162,EX163,EX164,EX165,EX166,EX167,EX168,EX169,EX170,
     EX171,EX172,EX173,EX174,EX175,EX176,EX177,EX178,EX179,EX180,
     EX181,EX182,EX183,EX184,EX185,EX186,EX187,EX188,EX189,EX190,
     EX191,EX192,EX193,EX194,EX195,EX196,EX197,EX198,EX199,EX200,
     EX201,EX202,EX203,EX204,EX205,EX206,EX207,EX208,EX209,EX210,
     EX211,EX212,EX213,EX214,EX215,EX216,EX217,EX218,EX219,EX220,
     EX221,EX222,EX223,EX224,EX225,EX226,EX227,EX228,EX229,EX230,
     EX231,EX232,EX233,EX234,EX235,EX236,EX237,EX238,EX239,EX240,
     EX241,EX242,EX243,EX244,EX245,EX246,EX247,EX248,EX249,EX250,
     EX251,EX252,EX253,EX254,EX255,EX256,EX257,EX258,EX259,EX260,
     EX261,EX262,EX263,EX264,EX265,EX266,EX267,EX268,EX269,EX270,
     EX271,EX272,EX273,EX274,EX275,EX276,EX277,EX278,EX279,EX280,
     EX281,EX282,EX283,EX284,EX285,EX286,EX287,EX288,EX289,EX290,
     EX291,EX292,EX293,EX294,EX295,EX296,EX297,EX298,EX299,EX300,
     EX301,EX302,EX303,EX304,EX305,EX306,EX307,EX308,EX309,EX310,
     EX311,EX312,EX313,EX314,EX315,EX316,EX317,EX318,EX319,EX320,
     EX321,EX322,EX323,EX324,EX325,EX326,EX327,EX328,EX329,EX330,
     EX331,EX332,EX333,EX334,EX335,EX336,EX337,EX338,EX339,EX340,
     EX341,EX342,EX343,EX344,EX345,EX346,EX347,EX348,EX349,EX350,
     EX351,EX352,EX353,EX354,EX355,EX356,EX357,EX358,EX359,EX360,
     EX361,EX362,EX363,EX364,EX365,EX366,EX367,EX368,EX369,EX370,
     EX371,EX372,EX373,EX374,EX375,EX376,EX377,EX378,EX379,EX380,
     EX381,EX382,EX383,EX384,EX385,EX386,EX387,EX388,EX389,EX390,
     EX391,EX392,EX393,EX394,EX395,EX396,EX397,EX398,EX399,EX400,
     EX401,EX402,EX403,EX404,EX405,EX406,EX407,EX408,EX409,EX410,
     EX411,EX412,EX413,EX414,EX415,EX416,EX417,EX418,EX419,EX420,
     EX421,EX422,EX423,EX424,EX425,EX426,EX427,EX428,EX429,EX430,
     EX431,EX432,EX433,EX434,EX435,EX436,EX437,EX438,EX439,EX440,
     EX441,EX442,EX443,EX444,EX445,EX446,EX447,EX448,EX449,EX450,
     EX451,EX452,EX453,EX454,EX455,EX456,EX457,EX458,EX459,EX460,
     EX461,EX462,EX463,EX464,EX465,EX466,EX467,EX468,EX469,EX470,
     EX471,EX472,EX473,EX474,EX475,EX476,EX477,EX478,EX479,EX480,
     EX481,EX482,EX483,EX484,EX485,EX486,EX487,EX488,EX489,EX490,
     EX491,EX492,EX493,EX494,EX495,EX496,EX497,EX498,EX499,EX500,
     EX501,EX502,EX503,EX504,EX505,EX506,EX507,EX508,EX509,EX510,
     EX511,EX512,EX513,EX514,EX515,EX516,EX517,EX518,EX519,EX520,
     EX521,EX522,EX523,EX524,EX525,EX526,EX527,EX528,EX529,EX530,
     EX531,EX532,EX533,EX534,EX535,EX536,EX537,EX538,EX539,EX540,
     EX541,EX542,EX543,EX544,EX545,EX546,EX547,EX548,EX549,EX550,
     EX551,EX552,EX553,EX554,EX555,EX556,EX557,EX558,EX559,EX560,
     EX561,EX562,EX563,EX564,EX565,EX566,EX567,EX568,EX569,EX570,
     EX571,EX572,EX573,EX574,EX575,EX576,EX577,EX578,EX579,EX580,
     EX581,EX582,EX583,EX584,EX585,EX586,EX587,EX588,EX589,EX590,
     EX591,EX592,EX593,EX594,EX595,EX596,EX597,EX598,EX599,EX600,
     EX601,EX602,EX603,EX604,EX605,EX606,EX607,EX608,EX609,EX610,
     EX611,EX612,EX613,EX614,EX615,EX616,EX617,EX618,EX619,EX620,
     EX621,EX622,EX623,EX624,EX625,EX626,EX627,EX628,EX629,EX630,
     EX631,EX632,EX633,EX634,EX635,EX636,EX637,EX638,EX639,EX640,
     EX641,EX642,EX643,EX644,EX645,EX646,EX647,EX648,EX649,EX650,
     EX651,EX652,EX653,EX654,EX655,EX656,EX657,EX658,EX659,EX660,
     EX661,EX662,EX663,EX664,EX665,EX666,EX667,EX668,EX669,EX670,
     EX671,EX672,EX673,EX674,EX675,EX676,EX677,EX678,EX679,EX680,
     EX681,EX682,EX683,EX684,EX685,EX686,EX687,EX688,EX689,EX690,
     EX691,EX692,EX693,EX694,EX695,EX696,EX697,EX698,EX699,EX700,
     EX701,EX702,EX703,EX704,EX705,EX706,EX707,EX708,EX709,EX710,
     EX711,EX712,EX713,EX714,EX715,EX716,EX717,EX718,EX719,EX720,
     EX721,EX722,EX723,EX724,EX725,EX726,EX727,EX728,EX729,EX730,
     EX731,EX732,EX733,EX734,EX735,EX736,EX737,EX738,EX739,EX740,
     EX741,EX742,EX743,EX744,EX745,EX746,EX747,EX748,EX749,EX750,
     EX751,EX752,EX753,EX754,EX755,EX756,EX757,EX758,EX759,EX760,
     EX761,EX762,EX763,EX764,EX765,EX766,EX767,EX768,EX769,EX770,
     EX771,EX772,EX773,EX774,EX775,EX776,EX777,EX778,EX779,EX780,
     EX781,EX782,EX783,EX784,EX785,EX786,EX787,EX788,EX789,EX790,
     EX791,EX792,EX793,EX794,EX795,EX796,EX797,EX798,EX799,EX800,
     EX801,EX802,EX803,EX804,EX805,EX806,EX807,EX808,EX809,EX810,
     EX811,EX812,EX813,EX814,EX815,EX816,EX817,EX818,EX819,EX820,
     EX821,EX822,EX823,EX824,EX825,EX826,EX827,EX828,EX829,EX830,
     EX831,EX832,EX833,EX834,EX835,EX836,EX837,EX838,EX839,EX840,
     EX841,EX842,EX843,EX844,EX845,EX846,EX847,EX848,EX849,EX850,
     EX851,EX852,EX853,EX854,EX855,EX856,EX857,EX858,EX859,EX860,
     EX861,EX862,EX863,EX864,EX865,EX866,EX867,EX868,EX869,EX870,
     EX871,EX872,EX873,EX874,EX875,EX876,EX877,EX878,EX879,EX880,
     EX881,EX882,EX883,EX884,EX885,EX886,EX887,EX888,EX889,EX890,
     EX891,EX892,EX893,EX894,EX895,EX896,EX897,EX898,EX899,EX900,
     EX901,EX902,EX903,EX904,EX905,EX906,EX907,EX908,EX909,EX910,
     EX911,EX912,EX913,EX914,EX915,EX916,EX917,EX918,EX919,EX920,
     EX921,EX922,EX923,EX924,EX925,EX926,EX927,EX928,EX929,EX930,
     EX931,EX932,EX933,EX934,EX935,EX936,EX937,EX938,EX939,EX940,
     EX941,EX942,EX943,EX944,EX945,EX946,EX947,EX948,EX949,EX950,
     EX951,EX952,EX953,EX954,EX955,EX956,EX957,EX958,EX959,EX960,
     EX961,EX962,EX963,EX964,EX965,EX966,EX967,EX968,EX969,EX970,
     EX971,EX972,EX973,EX974,EX975,EX976,EX977,EX978,EX979,EX980,
     EX981,EX982,EX983,EX984,EX985,EX986,EX987,EX988,EX989,EX990,
     EX991,EX992,EX993,EX994,EX995,EX996,EX997,EX998,EX999,EX1000,
     EX1001,EX1002,EX1003,EX1004,EX1005,EX1006,EX1007,EX1008,EX1009,EX1010,
     EX1011,EX1012,EX1013,EX1014,EX1015,EX1016,EX1017,EX1018,EX1019,EX1020,
     EX1021,EX1022,EX1023,EX1024,EX1025,EX1026,EX1027,EX1028,EX1029,EX1030,
     EX1031,EX1032,EX1033,EX1034,EX1035,EX1036,EX1037,EX1038,EX1039,EX1040,
     EX1041,EX1042,EX1043,EX1044,EX1045,EX1046,EX1047,EX1048,EX1049,EX1050,
     EX1051,EX1052,EX1053,EX1054,EX1055,EX1056,EX1057,EX1058,EX1059,EX1060,
     EX1061,EX1062,EX1063,EX1064,EX1065,EX1066,EX1067,EX1068,EX1069,EX1070,
     EX1071,EX1072,EX1073,EX1074,EX1075,EX1076,EX1077,EX1078,EX1079,EX1080,
     EX1081,EX1082,EX1083,EX1084,EX1085,EX1086,EX1087,EX1088,EX1089,EX1090,
     EX1091,EX1092,EX1093,EX1094,EX1095,EX1096,EX1097,EX1098,EX1099,EX1100,
     EX1101,EX1102,EX1103,EX1104,EX1105,EX1106,EX1107,EX1108,EX1109,EX1110;


nand4 gate1( .a(N1), .b(N8), .c(N13), .d(N17), .O(N269) );
nand4 gate2( .a(N1), .b(N26), .c(N13), .d(N17), .O(N270) );
and3 gate3( .a(N29), .b(N36), .c(N42), .O(N273) );
and3 gate4( .a(N1), .b(N26), .c(N51), .O(N276) );
nand4 gate5( .a(N1), .b(N8), .c(N51), .d(N17), .O(N279) );
nand4 gate6( .a(N1), .b(N8), .c(N13), .d(N55), .O(N280) );
nand4 gate7( .a(N59), .b(N42), .c(N68), .d(N72), .O(N284) );
nand2 gate8( .a(N29), .b(N68), .O(N285) );
nand3 gate9( .a(N59), .b(N68), .c(N74), .O(N286) );
and3 gate10( .a(N29), .b(N75), .c(N80), .O(N287) );
and3 gate11( .a(N29), .b(N75), .c(N42), .O(N290) );
and3 gate12( .a(N29), .b(N36), .c(N80), .O(N291) );
and3 gate13( .a(N29), .b(N36), .c(N42), .O(N292) );
and3 gate14( .a(N59), .b(N75), .c(N80), .O(N293) );
and3 gate15( .a(N59), .b(N75), .c(N42), .O(N294) );
and3 gate16( .a(N59), .b(N36), .c(N80), .O(N295) );
and3 gate17( .a(N59), .b(N36), .c(N42), .O(N296) );
and2 gate18( .a(N85), .b(N86), .O(N297) );
or2 gate19( .a(N87), .b(N88), .O(N298) );
nand2 gate20( .a(N91), .b(N96), .O(N301) );
or2 gate21( .a(N91), .b(N96), .O(N302) );
inv1 gate( .a(N101),.O(N101_NOT) );
inv1 gate( .a(N106),.O(N106_NOT));
and2 gate( .a(N101_NOT), .b(p1), .O(EX1) );
and2 gate( .a(N106_NOT), .b(EX1), .O(EX2) );
and2 gate( .a(N101), .b(p2), .O(EX3) );
and2 gate( .a(N106_NOT), .b(EX3), .O(EX4) );
and2 gate( .a(N101_NOT), .b(p3), .O(EX5) );
and2 gate( .a(N106), .b(EX5), .O(EX6) );
and2 gate( .a(N101), .b(p4), .O(EX7) );
and2 gate( .a(N106), .b(EX7), .O(EX8) );
or2  gate( .a(EX2), .b(EX4), .O(EX9) );
or2  gate( .a(EX6), .b(EX9), .O(EX10) );
or2  gate( .a(EX8), .b(EX10), .O(N303) );
inv1 gate( .a(N101),.O(N101_NOT) );
inv1 gate( .a(N106),.O(N106_NOT));
and2 gate( .a(N101_NOT), .b(p5), .O(EX11) );
and2 gate( .a(N106_NOT), .b(EX11), .O(EX12) );
and2 gate( .a(N101), .b(p6), .O(EX13) );
and2 gate( .a(N106_NOT), .b(EX13), .O(EX14) );
and2 gate( .a(N101_NOT), .b(p7), .O(EX15) );
and2 gate( .a(N106), .b(EX15), .O(EX16) );
and2 gate( .a(N101), .b(p8), .O(EX17) );
and2 gate( .a(N106), .b(EX17), .O(EX18) );
or2  gate( .a(EX12), .b(EX14), .O(EX19) );
or2  gate( .a(EX16), .b(EX19), .O(EX20) );
or2  gate( .a(EX18), .b(EX20), .O(N304) );
nand2 gate24( .a(N111), .b(N116), .O(N305) );
inv1 gate( .a(N111),.O(N111_NOT) );
inv1 gate( .a(N116),.O(N116_NOT));
and2 gate( .a(N111_NOT), .b(p9), .O(EX21) );
and2 gate( .a(N116_NOT), .b(EX21), .O(EX22) );
and2 gate( .a(N111), .b(p10), .O(EX23) );
and2 gate( .a(N116_NOT), .b(EX23), .O(EX24) );
and2 gate( .a(N111_NOT), .b(p11), .O(EX25) );
and2 gate( .a(N116), .b(EX25), .O(EX26) );
and2 gate( .a(N111), .b(p12), .O(EX27) );
and2 gate( .a(N116), .b(EX27), .O(EX28) );
or2  gate( .a(EX22), .b(EX24), .O(EX29) );
or2  gate( .a(EX26), .b(EX29), .O(EX30) );
or2  gate( .a(EX28), .b(EX30), .O(N306) );
inv1 gate( .a(N121),.O(N121_NOT) );
inv1 gate( .a(N126),.O(N126_NOT));
and2 gate( .a(N121_NOT), .b(p13), .O(EX31) );
and2 gate( .a(N126_NOT), .b(EX31), .O(EX32) );
and2 gate( .a(N121), .b(p14), .O(EX33) );
and2 gate( .a(N126_NOT), .b(EX33), .O(EX34) );
and2 gate( .a(N121_NOT), .b(p15), .O(EX35) );
and2 gate( .a(N126), .b(EX35), .O(EX36) );
and2 gate( .a(N121), .b(p16), .O(EX37) );
and2 gate( .a(N126), .b(EX37), .O(EX38) );
or2  gate( .a(EX32), .b(EX34), .O(EX39) );
or2  gate( .a(EX36), .b(EX39), .O(EX40) );
or2  gate( .a(EX38), .b(EX40), .O(N307) );
or2 gate27( .a(N121), .b(N126), .O(N308) );
and2 gate28( .a(N8), .b(N138), .O(N309) );
inv1 gate29( .a(N268), .O(N310) );
and2 gate30( .a(N51), .b(N138), .O(N316) );
inv1 gate( .a(N17),.O(N17_NOT) );
inv1 gate( .a(N138),.O(N138_NOT));
and2 gate( .a(N17_NOT), .b(p17), .O(EX41) );
and2 gate( .a(N138_NOT), .b(EX41), .O(EX42) );
and2 gate( .a(N17), .b(p18), .O(EX43) );
and2 gate( .a(N138_NOT), .b(EX43), .O(EX44) );
and2 gate( .a(N17_NOT), .b(p19), .O(EX45) );
and2 gate( .a(N138), .b(EX45), .O(EX46) );
and2 gate( .a(N17), .b(p20), .O(EX47) );
and2 gate( .a(N138), .b(EX47), .O(EX48) );
or2  gate( .a(EX42), .b(EX44), .O(EX49) );
or2  gate( .a(EX46), .b(EX49), .O(EX50) );
or2  gate( .a(EX48), .b(EX50), .O(N317) );
inv1 gate( .a(N152),.O(N152_NOT) );
inv1 gate( .a(N138),.O(N138_NOT));
and2 gate( .a(N152_NOT), .b(p21), .O(EX51) );
and2 gate( .a(N138_NOT), .b(EX51), .O(EX52) );
and2 gate( .a(N152), .b(p22), .O(EX53) );
and2 gate( .a(N138_NOT), .b(EX53), .O(EX54) );
and2 gate( .a(N152_NOT), .b(p23), .O(EX55) );
and2 gate( .a(N138), .b(EX55), .O(EX56) );
and2 gate( .a(N152), .b(p24), .O(EX57) );
and2 gate( .a(N138), .b(EX57), .O(EX58) );
or2  gate( .a(EX52), .b(EX54), .O(EX59) );
or2  gate( .a(EX56), .b(EX59), .O(EX60) );
or2  gate( .a(EX58), .b(EX60), .O(N318) );
nand2 gate33( .a(N59), .b(N156), .O(N319) );
nor2 gate34( .a(N17), .b(N42), .O(N322) );
inv1 gate( .a(N17),.O(N17_NOT) );
inv1 gate( .a(N42),.O(N42_NOT));
and2 gate( .a(N17_NOT), .b(p25), .O(EX61) );
and2 gate( .a(N42_NOT), .b(EX61), .O(EX62) );
and2 gate( .a(N17), .b(p26), .O(EX63) );
and2 gate( .a(N42_NOT), .b(EX63), .O(EX64) );
and2 gate( .a(N17_NOT), .b(p27), .O(EX65) );
and2 gate( .a(N42), .b(EX65), .O(EX66) );
and2 gate( .a(N17), .b(p28), .O(EX67) );
and2 gate( .a(N42), .b(EX67), .O(EX68) );
or2  gate( .a(EX62), .b(EX64), .O(EX69) );
or2  gate( .a(EX66), .b(EX69), .O(EX70) );
or2  gate( .a(EX68), .b(EX70), .O(N323) );
nand2 gate36( .a(N159), .b(N165), .O(N324) );
inv1 gate( .a(N159),.O(N159_NOT) );
inv1 gate( .a(N165),.O(N165_NOT));
and2 gate( .a(N159_NOT), .b(p29), .O(EX71) );
and2 gate( .a(N165_NOT), .b(EX71), .O(EX72) );
and2 gate( .a(N159), .b(p30), .O(EX73) );
and2 gate( .a(N165_NOT), .b(EX73), .O(EX74) );
and2 gate( .a(N159_NOT), .b(p31), .O(EX75) );
and2 gate( .a(N165), .b(EX75), .O(EX76) );
and2 gate( .a(N159), .b(p32), .O(EX77) );
and2 gate( .a(N165), .b(EX77), .O(EX78) );
or2  gate( .a(EX72), .b(EX74), .O(EX79) );
or2  gate( .a(EX76), .b(EX79), .O(EX80) );
or2  gate( .a(EX78), .b(EX80), .O(N325) );
inv1 gate( .a(N171),.O(N171_NOT) );
inv1 gate( .a(N177),.O(N177_NOT));
and2 gate( .a(N171_NOT), .b(p33), .O(EX81) );
and2 gate( .a(N177_NOT), .b(EX81), .O(EX82) );
and2 gate( .a(N171), .b(p34), .O(EX83) );
and2 gate( .a(N177_NOT), .b(EX83), .O(EX84) );
and2 gate( .a(N171_NOT), .b(p35), .O(EX85) );
and2 gate( .a(N177), .b(EX85), .O(EX86) );
and2 gate( .a(N171), .b(p36), .O(EX87) );
and2 gate( .a(N177), .b(EX87), .O(EX88) );
or2  gate( .a(EX82), .b(EX84), .O(EX89) );
or2  gate( .a(EX86), .b(EX89), .O(EX90) );
or2  gate( .a(EX88), .b(EX90), .O(N326) );
inv1 gate( .a(N171),.O(N171_NOT) );
inv1 gate( .a(N177),.O(N177_NOT));
and2 gate( .a(N171_NOT), .b(p37), .O(EX91) );
and2 gate( .a(N177_NOT), .b(EX91), .O(EX92) );
and2 gate( .a(N171), .b(p38), .O(EX93) );
and2 gate( .a(N177_NOT), .b(EX93), .O(EX94) );
and2 gate( .a(N171_NOT), .b(p39), .O(EX95) );
and2 gate( .a(N177), .b(EX95), .O(EX96) );
and2 gate( .a(N171), .b(p40), .O(EX97) );
and2 gate( .a(N177), .b(EX97), .O(EX98) );
or2  gate( .a(EX92), .b(EX94), .O(EX99) );
or2  gate( .a(EX96), .b(EX99), .O(EX100) );
or2  gate( .a(EX98), .b(EX100), .O(N327) );
nand2 gate40( .a(N183), .b(N189), .O(N328) );
or2 gate41( .a(N183), .b(N189), .O(N329) );
nand2 gate42( .a(N195), .b(N201), .O(N330) );
or2 gate43( .a(N195), .b(N201), .O(N331) );
and2 gate44( .a(N210), .b(N91), .O(N332) );
inv1 gate( .a(N210),.O(N210_NOT) );
inv1 gate( .a(N96),.O(N96_NOT));
and2 gate( .a(N210_NOT), .b(p41), .O(EX101) );
and2 gate( .a(N96_NOT), .b(EX101), .O(EX102) );
and2 gate( .a(N210), .b(p42), .O(EX103) );
and2 gate( .a(N96_NOT), .b(EX103), .O(EX104) );
and2 gate( .a(N210_NOT), .b(p43), .O(EX105) );
and2 gate( .a(N96), .b(EX105), .O(EX106) );
and2 gate( .a(N210), .b(p44), .O(EX107) );
and2 gate( .a(N96), .b(EX107), .O(EX108) );
or2  gate( .a(EX102), .b(EX104), .O(EX109) );
or2  gate( .a(EX106), .b(EX109), .O(EX110) );
or2  gate( .a(EX108), .b(EX110), .O(N333) );
and2 gate46( .a(N210), .b(N101), .O(N334) );
and2 gate47( .a(N210), .b(N106), .O(N335) );
inv1 gate( .a(N210),.O(N210_NOT) );
inv1 gate( .a(N111),.O(N111_NOT));
and2 gate( .a(N210_NOT), .b(p45), .O(EX111) );
and2 gate( .a(N111_NOT), .b(EX111), .O(EX112) );
and2 gate( .a(N210), .b(p46), .O(EX113) );
and2 gate( .a(N111_NOT), .b(EX113), .O(EX114) );
and2 gate( .a(N210_NOT), .b(p47), .O(EX115) );
and2 gate( .a(N111), .b(EX115), .O(EX116) );
and2 gate( .a(N210), .b(p48), .O(EX117) );
and2 gate( .a(N111), .b(EX117), .O(EX118) );
or2  gate( .a(EX112), .b(EX114), .O(EX119) );
or2  gate( .a(EX116), .b(EX119), .O(EX120) );
or2  gate( .a(EX118), .b(EX120), .O(N336) );
inv1 gate( .a(N255),.O(N255_NOT) );
inv1 gate( .a(N259),.O(N259_NOT));
and2 gate( .a(N255_NOT), .b(p49), .O(EX121) );
and2 gate( .a(N259_NOT), .b(EX121), .O(EX122) );
and2 gate( .a(N255), .b(p50), .O(EX123) );
and2 gate( .a(N259_NOT), .b(EX123), .O(EX124) );
and2 gate( .a(N255_NOT), .b(p51), .O(EX125) );
and2 gate( .a(N259), .b(EX125), .O(EX126) );
and2 gate( .a(N255), .b(p52), .O(EX127) );
and2 gate( .a(N259), .b(EX127), .O(EX128) );
or2  gate( .a(EX122), .b(EX124), .O(EX129) );
or2  gate( .a(EX126), .b(EX129), .O(EX130) );
or2  gate( .a(EX128), .b(EX130), .O(N337) );
inv1 gate( .a(N210),.O(N210_NOT) );
inv1 gate( .a(N116),.O(N116_NOT));
and2 gate( .a(N210_NOT), .b(p53), .O(EX131) );
and2 gate( .a(N116_NOT), .b(EX131), .O(EX132) );
and2 gate( .a(N210), .b(p54), .O(EX133) );
and2 gate( .a(N116_NOT), .b(EX133), .O(EX134) );
and2 gate( .a(N210_NOT), .b(p55), .O(EX135) );
and2 gate( .a(N116), .b(EX135), .O(EX136) );
and2 gate( .a(N210), .b(p56), .O(EX137) );
and2 gate( .a(N116), .b(EX137), .O(EX138) );
or2  gate( .a(EX132), .b(EX134), .O(EX139) );
or2  gate( .a(EX136), .b(EX139), .O(EX140) );
or2  gate( .a(EX138), .b(EX140), .O(N338) );
and2 gate51( .a(N255), .b(N260), .O(N339) );
and2 gate52( .a(N210), .b(N121), .O(N340) );
inv1 gate( .a(N255),.O(N255_NOT) );
inv1 gate( .a(N267),.O(N267_NOT));
and2 gate( .a(N255_NOT), .b(p57), .O(EX141) );
and2 gate( .a(N267_NOT), .b(EX141), .O(EX142) );
and2 gate( .a(N255), .b(p58), .O(EX143) );
and2 gate( .a(N267_NOT), .b(EX143), .O(EX144) );
and2 gate( .a(N255_NOT), .b(p59), .O(EX145) );
and2 gate( .a(N267), .b(EX145), .O(EX146) );
and2 gate( .a(N255), .b(p60), .O(EX147) );
and2 gate( .a(N267), .b(EX147), .O(EX148) );
or2  gate( .a(EX142), .b(EX144), .O(EX149) );
or2  gate( .a(EX146), .b(EX149), .O(EX150) );
or2  gate( .a(EX148), .b(EX150), .O(N341) );
inv1 gate54( .a(N269), .O(N342) );
inv1 gate55( .a(N273), .O(N343) );
inv1 gate( .a(N270),.O(N270_NOT) );
inv1 gate( .a(N273),.O(N273_NOT));
and2 gate( .a(N270_NOT), .b(p61), .O(EX151) );
and2 gate( .a(N273_NOT), .b(EX151), .O(EX152) );
and2 gate( .a(N270), .b(p62), .O(EX153) );
and2 gate( .a(N273_NOT), .b(EX153), .O(EX154) );
and2 gate( .a(N270_NOT), .b(p63), .O(EX155) );
and2 gate( .a(N273), .b(EX155), .O(EX156) );
and2 gate( .a(N270), .b(p64), .O(EX157) );
and2 gate( .a(N273), .b(EX157), .O(EX158) );
or2  gate( .a(EX152), .b(EX154), .O(EX159) );
or2  gate( .a(EX156), .b(EX159), .O(EX160) );
or2  gate( .a(EX158), .b(EX160), .O(N344) );
inv1 gate57( .a(N276), .O(N345) );
inv1 gate58( .a(N276), .O(N346) );
inv1 gate59( .a(N279), .O(N347) );
nor2 gate60( .a(N280), .b(N284), .O(N348) );
or2 gate61( .a(N280), .b(N285), .O(N349) );
inv1 gate( .a(N280),.O(N280_NOT) );
inv1 gate( .a(N286),.O(N286_NOT));
and2 gate( .a(N280_NOT), .b(p65), .O(EX161) );
and2 gate( .a(N286_NOT), .b(EX161), .O(EX162) );
and2 gate( .a(N280), .b(p66), .O(EX163) );
and2 gate( .a(N286_NOT), .b(EX163), .O(EX164) );
and2 gate( .a(N280_NOT), .b(p67), .O(EX165) );
and2 gate( .a(N286), .b(EX165), .O(EX166) );
and2 gate( .a(N280), .b(p68), .O(EX167) );
and2 gate( .a(N286), .b(EX167), .O(EX168) );
or2  gate( .a(EX162), .b(EX164), .O(EX169) );
or2  gate( .a(EX166), .b(EX169), .O(EX170) );
or2  gate( .a(EX168), .b(EX170), .O(N350) );
inv1 gate63( .a(N293), .O(N351) );
inv1 gate64( .a(N294), .O(N352) );
inv1 gate65( .a(N295), .O(N353) );
inv1 gate66( .a(N296), .O(N354) );
nand2 gate67( .a(N89), .b(N298), .O(N355) );
and2 gate68( .a(N90), .b(N298), .O(N356) );
nand2 gate69( .a(N301), .b(N302), .O(N357) );
nand2 gate70( .a(N303), .b(N304), .O(N360) );
inv1 gate( .a(N305),.O(N305_NOT) );
inv1 gate( .a(N306),.O(N306_NOT));
and2 gate( .a(N305_NOT), .b(p69), .O(EX171) );
and2 gate( .a(N306_NOT), .b(EX171), .O(EX172) );
and2 gate( .a(N305), .b(p70), .O(EX173) );
and2 gate( .a(N306_NOT), .b(EX173), .O(EX174) );
and2 gate( .a(N305_NOT), .b(p71), .O(EX175) );
and2 gate( .a(N306), .b(EX175), .O(EX176) );
and2 gate( .a(N305), .b(p72), .O(EX177) );
and2 gate( .a(N306), .b(EX177), .O(EX178) );
or2  gate( .a(EX172), .b(EX174), .O(EX179) );
or2  gate( .a(EX176), .b(EX179), .O(EX180) );
or2  gate( .a(EX178), .b(EX180), .O(N363) );
inv1 gate( .a(N307),.O(N307_NOT) );
inv1 gate( .a(N308),.O(N308_NOT));
and2 gate( .a(N307_NOT), .b(p73), .O(EX181) );
and2 gate( .a(N308_NOT), .b(EX181), .O(EX182) );
and2 gate( .a(N307), .b(p74), .O(EX183) );
and2 gate( .a(N308_NOT), .b(EX183), .O(EX184) );
and2 gate( .a(N307_NOT), .b(p75), .O(EX185) );
and2 gate( .a(N308), .b(EX185), .O(EX186) );
and2 gate( .a(N307), .b(p76), .O(EX187) );
and2 gate( .a(N308), .b(EX187), .O(EX188) );
or2  gate( .a(EX182), .b(EX184), .O(EX189) );
or2  gate( .a(EX186), .b(EX189), .O(EX190) );
or2  gate( .a(EX188), .b(EX190), .O(N366) );
inv1 gate73( .a(N310), .O(N369) );
inv1 gate( .a(N322),.O(N322_NOT) );
inv1 gate( .a(N323),.O(N323_NOT));
and2 gate( .a(N322_NOT), .b(p77), .O(EX191) );
and2 gate( .a(N323_NOT), .b(EX191), .O(EX192) );
and2 gate( .a(N322), .b(p78), .O(EX193) );
and2 gate( .a(N323_NOT), .b(EX193), .O(EX194) );
and2 gate( .a(N322_NOT), .b(p79), .O(EX195) );
and2 gate( .a(N323), .b(EX195), .O(EX196) );
and2 gate( .a(N322), .b(p80), .O(EX197) );
and2 gate( .a(N323), .b(EX197), .O(EX198) );
or2  gate( .a(EX192), .b(EX194), .O(EX199) );
or2  gate( .a(EX196), .b(EX199), .O(EX200) );
or2  gate( .a(EX198), .b(EX200), .O(N375) );
nand2 gate75( .a(N324), .b(N325), .O(N376) );
inv1 gate( .a(N326),.O(N326_NOT) );
inv1 gate( .a(N327),.O(N327_NOT));
and2 gate( .a(N326_NOT), .b(p81), .O(EX201) );
and2 gate( .a(N327_NOT), .b(EX201), .O(EX202) );
and2 gate( .a(N326), .b(p82), .O(EX203) );
and2 gate( .a(N327_NOT), .b(EX203), .O(EX204) );
and2 gate( .a(N326_NOT), .b(p83), .O(EX205) );
and2 gate( .a(N327), .b(EX205), .O(EX206) );
and2 gate( .a(N326), .b(p84), .O(EX207) );
and2 gate( .a(N327), .b(EX207), .O(EX208) );
or2  gate( .a(EX202), .b(EX204), .O(EX209) );
or2  gate( .a(EX206), .b(EX209), .O(EX210) );
or2  gate( .a(EX208), .b(EX210), .O(N379) );
nand2 gate77( .a(N328), .b(N329), .O(N382) );
inv1 gate( .a(N330),.O(N330_NOT) );
inv1 gate( .a(N331),.O(N331_NOT));
and2 gate( .a(N330_NOT), .b(p85), .O(EX211) );
and2 gate( .a(N331_NOT), .b(EX211), .O(EX212) );
and2 gate( .a(N330), .b(p86), .O(EX213) );
and2 gate( .a(N331_NOT), .b(EX213), .O(EX214) );
and2 gate( .a(N330_NOT), .b(p87), .O(EX215) );
and2 gate( .a(N331), .b(EX215), .O(EX216) );
and2 gate( .a(N330), .b(p88), .O(EX217) );
and2 gate( .a(N331), .b(EX217), .O(EX218) );
or2  gate( .a(EX212), .b(EX214), .O(EX219) );
or2  gate( .a(EX216), .b(EX219), .O(EX220) );
or2  gate( .a(EX218), .b(EX220), .O(N385) );
buf1 gate79( .a(N290), .O(N388) );
buf1 gate80( .a(N291), .O(N389) );
buf1 gate81( .a(N292), .O(N390) );
buf1 gate82( .a(N297), .O(N391) );
or2 gate83( .a(N270), .b(N343), .O(N392) );
inv1 gate84( .a(N345), .O(N393) );
inv1 gate85( .a(N346), .O(N399) );
inv1 gate( .a(N348),.O(N348_NOT) );
inv1 gate( .a(N73),.O(N73_NOT));
and2 gate( .a(N348_NOT), .b(p89), .O(EX221) );
and2 gate( .a(N73_NOT), .b(EX221), .O(EX222) );
and2 gate( .a(N348), .b(p90), .O(EX223) );
and2 gate( .a(N73_NOT), .b(EX223), .O(EX224) );
and2 gate( .a(N348_NOT), .b(p91), .O(EX225) );
and2 gate( .a(N73), .b(EX225), .O(EX226) );
and2 gate( .a(N348), .b(p92), .O(EX227) );
and2 gate( .a(N73), .b(EX227), .O(EX228) );
or2  gate( .a(EX222), .b(EX224), .O(EX229) );
or2  gate( .a(EX226), .b(EX229), .O(EX230) );
or2  gate( .a(EX228), .b(EX230), .O(N400) );
inv1 gate87( .a(N349), .O(N401) );
inv1 gate88( .a(N350), .O(N402) );
inv1 gate89( .a(N355), .O(N403) );
inv1 gate90( .a(N357), .O(N404) );
inv1 gate91( .a(N360), .O(N405) );
inv1 gate( .a(N357),.O(N357_NOT) );
inv1 gate( .a(N360),.O(N360_NOT));
and2 gate( .a(N357_NOT), .b(p93), .O(EX231) );
and2 gate( .a(N360_NOT), .b(EX231), .O(EX232) );
and2 gate( .a(N357), .b(p94), .O(EX233) );
and2 gate( .a(N360_NOT), .b(EX233), .O(EX234) );
and2 gate( .a(N357_NOT), .b(p95), .O(EX235) );
and2 gate( .a(N360), .b(EX235), .O(EX236) );
and2 gate( .a(N357), .b(p96), .O(EX237) );
and2 gate( .a(N360), .b(EX237), .O(EX238) );
or2  gate( .a(EX232), .b(EX234), .O(EX239) );
or2  gate( .a(EX236), .b(EX239), .O(EX240) );
or2  gate( .a(EX238), .b(EX240), .O(N406) );
inv1 gate93( .a(N363), .O(N407) );
inv1 gate94( .a(N366), .O(N408) );
inv1 gate( .a(N363),.O(N363_NOT) );
inv1 gate( .a(N366),.O(N366_NOT));
and2 gate( .a(N363_NOT), .b(p97), .O(EX241) );
and2 gate( .a(N366_NOT), .b(EX241), .O(EX242) );
and2 gate( .a(N363), .b(p98), .O(EX243) );
and2 gate( .a(N366_NOT), .b(EX243), .O(EX244) );
and2 gate( .a(N363_NOT), .b(p99), .O(EX245) );
and2 gate( .a(N366), .b(EX245), .O(EX246) );
and2 gate( .a(N363), .b(p100), .O(EX247) );
and2 gate( .a(N366), .b(EX247), .O(EX248) );
or2  gate( .a(EX242), .b(EX244), .O(EX249) );
or2  gate( .a(EX246), .b(EX249), .O(EX250) );
or2  gate( .a(EX248), .b(EX250), .O(N409) );
nand2 gate96( .a(N347), .b(N352), .O(N410) );
inv1 gate97( .a(N376), .O(N411) );
inv1 gate98( .a(N379), .O(N412) );
and2 gate99( .a(N376), .b(N379), .O(N413) );
inv1 gate100( .a(N382), .O(N414) );
inv1 gate101( .a(N385), .O(N415) );
and2 gate102( .a(N382), .b(N385), .O(N416) );
inv1 gate( .a(N210),.O(N210_NOT) );
inv1 gate( .a(N369),.O(N369_NOT));
and2 gate( .a(N210_NOT), .b(p101), .O(EX251) );
and2 gate( .a(N369_NOT), .b(EX251), .O(EX252) );
and2 gate( .a(N210), .b(p102), .O(EX253) );
and2 gate( .a(N369_NOT), .b(EX253), .O(EX254) );
and2 gate( .a(N210_NOT), .b(p103), .O(EX255) );
and2 gate( .a(N369), .b(EX255), .O(EX256) );
and2 gate( .a(N210), .b(p104), .O(EX257) );
and2 gate( .a(N369), .b(EX257), .O(EX258) );
or2  gate( .a(EX252), .b(EX254), .O(EX259) );
or2  gate( .a(EX256), .b(EX259), .O(EX260) );
or2  gate( .a(EX258), .b(EX260), .O(N417) );
buf1 gate104( .a(N342), .O(N418) );
buf1 gate105( .a(N344), .O(N419) );
buf1 gate106( .a(N351), .O(N420) );
buf1 gate107( .a(N353), .O(N421) );
buf1 gate108( .a(N354), .O(N422) );
buf1 gate109( .a(N356), .O(N423) );
inv1 gate110( .a(N400), .O(N424) );
and2 gate111( .a(N404), .b(N405), .O(N425) );
inv1 gate( .a(N407),.O(N407_NOT) );
inv1 gate( .a(N408),.O(N408_NOT));
and2 gate( .a(N407_NOT), .b(p105), .O(EX261) );
and2 gate( .a(N408_NOT), .b(EX261), .O(EX262) );
and2 gate( .a(N407), .b(p106), .O(EX263) );
and2 gate( .a(N408_NOT), .b(EX263), .O(EX264) );
and2 gate( .a(N407_NOT), .b(p107), .O(EX265) );
and2 gate( .a(N408), .b(EX265), .O(EX266) );
and2 gate( .a(N407), .b(p108), .O(EX267) );
and2 gate( .a(N408), .b(EX267), .O(EX268) );
or2  gate( .a(EX262), .b(EX264), .O(EX269) );
or2  gate( .a(EX266), .b(EX269), .O(EX270) );
or2  gate( .a(EX268), .b(EX270), .O(N426) );
and3 gate113( .a(N319), .b(N393), .c(N55), .O(N427) );
and3 gate114( .a(N393), .b(N17), .c(N287), .O(N432) );
nand3 gate115( .a(N393), .b(N287), .c(N55), .O(N437) );
nand4 gate116( .a(N375), .b(N59), .c(N156), .d(N393), .O(N442) );
nand3 gate117( .a(N393), .b(N319), .c(N17), .O(N443) );
inv1 gate( .a(N411),.O(N411_NOT) );
inv1 gate( .a(N412),.O(N412_NOT));
and2 gate( .a(N411_NOT), .b(p109), .O(EX271) );
and2 gate( .a(N412_NOT), .b(EX271), .O(EX272) );
and2 gate( .a(N411), .b(p110), .O(EX273) );
and2 gate( .a(N412_NOT), .b(EX273), .O(EX274) );
and2 gate( .a(N411_NOT), .b(p111), .O(EX275) );
and2 gate( .a(N412), .b(EX275), .O(EX276) );
and2 gate( .a(N411), .b(p112), .O(EX277) );
and2 gate( .a(N412), .b(EX277), .O(EX278) );
or2  gate( .a(EX272), .b(EX274), .O(EX279) );
or2  gate( .a(EX276), .b(EX279), .O(EX280) );
or2  gate( .a(EX278), .b(EX280), .O(N444) );
and2 gate119( .a(N414), .b(N415), .O(N445) );
buf1 gate120( .a(N392), .O(N446) );
buf1 gate121( .a(N399), .O(N447) );
buf1 gate122( .a(N401), .O(N448) );
buf1 gate123( .a(N402), .O(N449) );
buf1 gate124( .a(N403), .O(N450) );
inv1 gate125( .a(N424), .O(N451) );
nor2 gate126( .a(N406), .b(N425), .O(N460) );
nor2 gate127( .a(N409), .b(N426), .O(N463) );
inv1 gate( .a(N442),.O(N442_NOT) );
inv1 gate( .a(N410),.O(N410_NOT));
and2 gate( .a(N442_NOT), .b(p113), .O(EX281) );
and2 gate( .a(N410_NOT), .b(EX281), .O(EX282) );
and2 gate( .a(N442), .b(p114), .O(EX283) );
and2 gate( .a(N410_NOT), .b(EX283), .O(EX284) );
and2 gate( .a(N442_NOT), .b(p115), .O(EX285) );
and2 gate( .a(N410), .b(EX285), .O(EX286) );
and2 gate( .a(N442), .b(p116), .O(EX287) );
and2 gate( .a(N410), .b(EX287), .O(EX288) );
or2  gate( .a(EX282), .b(EX284), .O(EX289) );
or2  gate( .a(EX286), .b(EX289), .O(EX290) );
or2  gate( .a(EX288), .b(EX290), .O(N466) );
inv1 gate( .a(N143),.O(N143_NOT) );
inv1 gate( .a(N427),.O(N427_NOT));
and2 gate( .a(N143_NOT), .b(p117), .O(EX291) );
and2 gate( .a(N427_NOT), .b(EX291), .O(EX292) );
and2 gate( .a(N143), .b(p118), .O(EX293) );
and2 gate( .a(N427_NOT), .b(EX293), .O(EX294) );
and2 gate( .a(N143_NOT), .b(p119), .O(EX295) );
and2 gate( .a(N427), .b(EX295), .O(EX296) );
and2 gate( .a(N143), .b(p120), .O(EX297) );
and2 gate( .a(N427), .b(EX297), .O(EX298) );
or2  gate( .a(EX292), .b(EX294), .O(EX299) );
or2  gate( .a(EX296), .b(EX299), .O(EX300) );
or2  gate( .a(EX298), .b(EX300), .O(N475) );
and2 gate130( .a(N310), .b(N432), .O(N476) );
and2 gate131( .a(N146), .b(N427), .O(N477) );
and2 gate132( .a(N310), .b(N432), .O(N478) );
and2 gate133( .a(N149), .b(N427), .O(N479) );
inv1 gate( .a(N310),.O(N310_NOT) );
inv1 gate( .a(N432),.O(N432_NOT));
and2 gate( .a(N310_NOT), .b(p121), .O(EX301) );
and2 gate( .a(N432_NOT), .b(EX301), .O(EX302) );
and2 gate( .a(N310), .b(p122), .O(EX303) );
and2 gate( .a(N432_NOT), .b(EX303), .O(EX304) );
and2 gate( .a(N310_NOT), .b(p123), .O(EX305) );
and2 gate( .a(N432), .b(EX305), .O(EX306) );
and2 gate( .a(N310), .b(p124), .O(EX307) );
and2 gate( .a(N432), .b(EX307), .O(EX308) );
or2  gate( .a(EX302), .b(EX304), .O(EX309) );
or2  gate( .a(EX306), .b(EX309), .O(EX310) );
or2  gate( .a(EX308), .b(EX310), .O(N480) );
and2 gate135( .a(N153), .b(N427), .O(N481) );
and2 gate136( .a(N310), .b(N432), .O(N482) );
inv1 gate( .a(N443),.O(N443_NOT) );
inv1 gate( .a(N1),.O(N1_NOT));
and2 gate( .a(N443_NOT), .b(p125), .O(EX311) );
and2 gate( .a(N1_NOT), .b(EX311), .O(EX312) );
and2 gate( .a(N443), .b(p126), .O(EX313) );
and2 gate( .a(N1_NOT), .b(EX313), .O(EX314) );
and2 gate( .a(N443_NOT), .b(p127), .O(EX315) );
and2 gate( .a(N1), .b(EX315), .O(EX316) );
and2 gate( .a(N443), .b(p128), .O(EX317) );
and2 gate( .a(N1), .b(EX317), .O(EX318) );
or2  gate( .a(EX312), .b(EX314), .O(EX319) );
or2  gate( .a(EX316), .b(EX319), .O(EX320) );
or2  gate( .a(EX318), .b(EX320), .O(N483) );
or2 gate138( .a(N369), .b(N437), .O(N488) );
inv1 gate( .a(N369),.O(N369_NOT) );
inv1 gate( .a(N437),.O(N437_NOT));
and2 gate( .a(N369_NOT), .b(p129), .O(EX321) );
and2 gate( .a(N437_NOT), .b(EX321), .O(EX322) );
and2 gate( .a(N369), .b(p130), .O(EX323) );
and2 gate( .a(N437_NOT), .b(EX323), .O(EX324) );
and2 gate( .a(N369_NOT), .b(p131), .O(EX325) );
and2 gate( .a(N437), .b(EX325), .O(EX326) );
and2 gate( .a(N369), .b(p132), .O(EX327) );
and2 gate( .a(N437), .b(EX327), .O(EX328) );
or2  gate( .a(EX322), .b(EX324), .O(EX329) );
or2  gate( .a(EX326), .b(EX329), .O(EX330) );
or2  gate( .a(EX328), .b(EX330), .O(N489) );
or2 gate140( .a(N369), .b(N437), .O(N490) );
or2 gate141( .a(N369), .b(N437), .O(N491) );
nor2 gate142( .a(N413), .b(N444), .O(N492) );
nor2 gate143( .a(N416), .b(N445), .O(N495) );
inv1 gate( .a(N130),.O(N130_NOT) );
inv1 gate( .a(N460),.O(N460_NOT));
and2 gate( .a(N130_NOT), .b(p133), .O(EX331) );
and2 gate( .a(N460_NOT), .b(EX331), .O(EX332) );
and2 gate( .a(N130), .b(p134), .O(EX333) );
and2 gate( .a(N460_NOT), .b(EX333), .O(EX334) );
and2 gate( .a(N130_NOT), .b(p135), .O(EX335) );
and2 gate( .a(N460), .b(EX335), .O(EX336) );
and2 gate( .a(N130), .b(p136), .O(EX337) );
and2 gate( .a(N460), .b(EX337), .O(EX338) );
or2  gate( .a(EX332), .b(EX334), .O(EX339) );
or2  gate( .a(EX336), .b(EX339), .O(EX340) );
or2  gate( .a(EX338), .b(EX340), .O(N498) );
inv1 gate( .a(N130),.O(N130_NOT) );
inv1 gate( .a(N460),.O(N460_NOT));
and2 gate( .a(N130_NOT), .b(p137), .O(EX341) );
and2 gate( .a(N460_NOT), .b(EX341), .O(EX342) );
and2 gate( .a(N130), .b(p138), .O(EX343) );
and2 gate( .a(N460_NOT), .b(EX343), .O(EX344) );
and2 gate( .a(N130_NOT), .b(p139), .O(EX345) );
and2 gate( .a(N460), .b(EX345), .O(EX346) );
and2 gate( .a(N130), .b(p140), .O(EX347) );
and2 gate( .a(N460), .b(EX347), .O(EX348) );
or2  gate( .a(EX342), .b(EX344), .O(EX349) );
or2  gate( .a(EX346), .b(EX349), .O(EX350) );
or2  gate( .a(EX348), .b(EX350), .O(N499) );
inv1 gate( .a(N463),.O(N463_NOT) );
inv1 gate( .a(N135),.O(N135_NOT));
and2 gate( .a(N463_NOT), .b(p141), .O(EX351) );
and2 gate( .a(N135_NOT), .b(EX351), .O(EX352) );
and2 gate( .a(N463), .b(p142), .O(EX353) );
and2 gate( .a(N135_NOT), .b(EX353), .O(EX354) );
and2 gate( .a(N463_NOT), .b(p143), .O(EX355) );
and2 gate( .a(N135), .b(EX355), .O(EX356) );
and2 gate( .a(N463), .b(p144), .O(EX357) );
and2 gate( .a(N135), .b(EX357), .O(EX358) );
or2  gate( .a(EX352), .b(EX354), .O(EX359) );
or2  gate( .a(EX356), .b(EX359), .O(EX360) );
or2  gate( .a(EX358), .b(EX360), .O(N500) );
or2 gate147( .a(N463), .b(N135), .O(N501) );
inv1 gate( .a(N91),.O(N91_NOT) );
inv1 gate( .a(N466),.O(N466_NOT));
and2 gate( .a(N91_NOT), .b(p145), .O(EX361) );
and2 gate( .a(N466_NOT), .b(EX361), .O(EX362) );
and2 gate( .a(N91), .b(p146), .O(EX363) );
and2 gate( .a(N466_NOT), .b(EX363), .O(EX364) );
and2 gate( .a(N91_NOT), .b(p147), .O(EX365) );
and2 gate( .a(N466), .b(EX365), .O(EX366) );
and2 gate( .a(N91), .b(p148), .O(EX367) );
and2 gate( .a(N466), .b(EX367), .O(EX368) );
or2  gate( .a(EX362), .b(EX364), .O(EX369) );
or2  gate( .a(EX366), .b(EX369), .O(EX370) );
or2  gate( .a(EX368), .b(EX370), .O(N502) );
inv1 gate( .a(N475),.O(N475_NOT) );
inv1 gate( .a(N476),.O(N476_NOT));
and2 gate( .a(N475_NOT), .b(p149), .O(EX371) );
and2 gate( .a(N476_NOT), .b(EX371), .O(EX372) );
and2 gate( .a(N475), .b(p150), .O(EX373) );
and2 gate( .a(N476_NOT), .b(EX373), .O(EX374) );
and2 gate( .a(N475_NOT), .b(p151), .O(EX375) );
and2 gate( .a(N476), .b(EX375), .O(EX376) );
and2 gate( .a(N475), .b(p152), .O(EX377) );
and2 gate( .a(N476), .b(EX377), .O(EX378) );
or2  gate( .a(EX372), .b(EX374), .O(EX379) );
or2  gate( .a(EX376), .b(EX379), .O(EX380) );
or2  gate( .a(EX378), .b(EX380), .O(N503) );
inv1 gate( .a(N96),.O(N96_NOT) );
inv1 gate( .a(N466),.O(N466_NOT));
and2 gate( .a(N96_NOT), .b(p153), .O(EX381) );
and2 gate( .a(N466_NOT), .b(EX381), .O(EX382) );
and2 gate( .a(N96), .b(p154), .O(EX383) );
and2 gate( .a(N466_NOT), .b(EX383), .O(EX384) );
and2 gate( .a(N96_NOT), .b(p155), .O(EX385) );
and2 gate( .a(N466), .b(EX385), .O(EX386) );
and2 gate( .a(N96), .b(p156), .O(EX387) );
and2 gate( .a(N466), .b(EX387), .O(EX388) );
or2  gate( .a(EX382), .b(EX384), .O(EX389) );
or2  gate( .a(EX386), .b(EX389), .O(EX390) );
or2  gate( .a(EX388), .b(EX390), .O(N504) );
inv1 gate( .a(N477),.O(N477_NOT) );
inv1 gate( .a(N478),.O(N478_NOT));
and2 gate( .a(N477_NOT), .b(p157), .O(EX391) );
and2 gate( .a(N478_NOT), .b(EX391), .O(EX392) );
and2 gate( .a(N477), .b(p158), .O(EX393) );
and2 gate( .a(N478_NOT), .b(EX393), .O(EX394) );
and2 gate( .a(N477_NOT), .b(p159), .O(EX395) );
and2 gate( .a(N478), .b(EX395), .O(EX396) );
and2 gate( .a(N477), .b(p160), .O(EX397) );
and2 gate( .a(N478), .b(EX397), .O(EX398) );
or2  gate( .a(EX392), .b(EX394), .O(EX399) );
or2  gate( .a(EX396), .b(EX399), .O(EX400) );
or2  gate( .a(EX398), .b(EX400), .O(N505) );
inv1 gate( .a(N101),.O(N101_NOT) );
inv1 gate( .a(N466),.O(N466_NOT));
and2 gate( .a(N101_NOT), .b(p161), .O(EX401) );
and2 gate( .a(N466_NOT), .b(EX401), .O(EX402) );
and2 gate( .a(N101), .b(p162), .O(EX403) );
and2 gate( .a(N466_NOT), .b(EX403), .O(EX404) );
and2 gate( .a(N101_NOT), .b(p163), .O(EX405) );
and2 gate( .a(N466), .b(EX405), .O(EX406) );
and2 gate( .a(N101), .b(p164), .O(EX407) );
and2 gate( .a(N466), .b(EX407), .O(EX408) );
or2  gate( .a(EX402), .b(EX404), .O(EX409) );
or2  gate( .a(EX406), .b(EX409), .O(EX410) );
or2  gate( .a(EX408), .b(EX410), .O(N506) );
nor2 gate153( .a(N479), .b(N480), .O(N507) );
and2 gate154( .a(N106), .b(N466), .O(N508) );
nor2 gate155( .a(N481), .b(N482), .O(N509) );
and2 gate156( .a(N143), .b(N483), .O(N510) );
and2 gate157( .a(N111), .b(N466), .O(N511) );
inv1 gate( .a(N146),.O(N146_NOT) );
inv1 gate( .a(N483),.O(N483_NOT));
and2 gate( .a(N146_NOT), .b(p165), .O(EX411) );
and2 gate( .a(N483_NOT), .b(EX411), .O(EX412) );
and2 gate( .a(N146), .b(p166), .O(EX413) );
and2 gate( .a(N483_NOT), .b(EX413), .O(EX414) );
and2 gate( .a(N146_NOT), .b(p167), .O(EX415) );
and2 gate( .a(N483), .b(EX415), .O(EX416) );
and2 gate( .a(N146), .b(p168), .O(EX417) );
and2 gate( .a(N483), .b(EX417), .O(EX418) );
or2  gate( .a(EX412), .b(EX414), .O(EX419) );
or2  gate( .a(EX416), .b(EX419), .O(EX420) );
or2  gate( .a(EX418), .b(EX420), .O(N512) );
inv1 gate( .a(N116),.O(N116_NOT) );
inv1 gate( .a(N466),.O(N466_NOT));
and2 gate( .a(N116_NOT), .b(p169), .O(EX421) );
and2 gate( .a(N466_NOT), .b(EX421), .O(EX422) );
and2 gate( .a(N116), .b(p170), .O(EX423) );
and2 gate( .a(N466_NOT), .b(EX423), .O(EX424) );
and2 gate( .a(N116_NOT), .b(p171), .O(EX425) );
and2 gate( .a(N466), .b(EX425), .O(EX426) );
and2 gate( .a(N116), .b(p172), .O(EX427) );
and2 gate( .a(N466), .b(EX427), .O(EX428) );
or2  gate( .a(EX422), .b(EX424), .O(EX429) );
or2  gate( .a(EX426), .b(EX429), .O(EX430) );
or2  gate( .a(EX428), .b(EX430), .O(N513) );
and2 gate160( .a(N149), .b(N483), .O(N514) );
and2 gate161( .a(N121), .b(N466), .O(N515) );
inv1 gate( .a(N153),.O(N153_NOT) );
inv1 gate( .a(N483),.O(N483_NOT));
and2 gate( .a(N153_NOT), .b(p173), .O(EX431) );
and2 gate( .a(N483_NOT), .b(EX431), .O(EX432) );
and2 gate( .a(N153), .b(p174), .O(EX433) );
and2 gate( .a(N483_NOT), .b(EX433), .O(EX434) );
and2 gate( .a(N153_NOT), .b(p175), .O(EX435) );
and2 gate( .a(N483), .b(EX435), .O(EX436) );
and2 gate( .a(N153), .b(p176), .O(EX437) );
and2 gate( .a(N483), .b(EX437), .O(EX438) );
or2  gate( .a(EX432), .b(EX434), .O(EX439) );
or2  gate( .a(EX436), .b(EX439), .O(EX440) );
or2  gate( .a(EX438), .b(EX440), .O(N516) );
and2 gate163( .a(N126), .b(N466), .O(N517) );
nand2 gate164( .a(N130), .b(N492), .O(N518) );
inv1 gate( .a(N130),.O(N130_NOT) );
inv1 gate( .a(N492),.O(N492_NOT));
and2 gate( .a(N130_NOT), .b(p177), .O(EX441) );
and2 gate( .a(N492_NOT), .b(EX441), .O(EX442) );
and2 gate( .a(N130), .b(p178), .O(EX443) );
and2 gate( .a(N492_NOT), .b(EX443), .O(EX444) );
and2 gate( .a(N130_NOT), .b(p179), .O(EX445) );
and2 gate( .a(N492), .b(EX445), .O(EX446) );
and2 gate( .a(N130), .b(p180), .O(EX447) );
and2 gate( .a(N492), .b(EX447), .O(EX448) );
or2  gate( .a(EX442), .b(EX444), .O(EX449) );
or2  gate( .a(EX446), .b(EX449), .O(EX450) );
or2  gate( .a(EX448), .b(EX450), .O(N519) );
nand2 gate166( .a(N495), .b(N207), .O(N520) );
inv1 gate( .a(N495),.O(N495_NOT) );
inv1 gate( .a(N207),.O(N207_NOT));
and2 gate( .a(N495_NOT), .b(p181), .O(EX451) );
and2 gate( .a(N207_NOT), .b(EX451), .O(EX452) );
and2 gate( .a(N495), .b(p182), .O(EX453) );
and2 gate( .a(N207_NOT), .b(EX453), .O(EX454) );
and2 gate( .a(N495_NOT), .b(p183), .O(EX455) );
and2 gate( .a(N207), .b(EX455), .O(EX456) );
and2 gate( .a(N495), .b(p184), .O(EX457) );
and2 gate( .a(N207), .b(EX457), .O(EX458) );
or2  gate( .a(EX452), .b(EX454), .O(EX459) );
or2  gate( .a(EX456), .b(EX459), .O(EX460) );
or2  gate( .a(EX458), .b(EX460), .O(N521) );
and2 gate168( .a(N451), .b(N159), .O(N522) );
inv1 gate( .a(N451),.O(N451_NOT) );
inv1 gate( .a(N165),.O(N165_NOT));
and2 gate( .a(N451_NOT), .b(p185), .O(EX461) );
and2 gate( .a(N165_NOT), .b(EX461), .O(EX462) );
and2 gate( .a(N451), .b(p186), .O(EX463) );
and2 gate( .a(N165_NOT), .b(EX463), .O(EX464) );
and2 gate( .a(N451_NOT), .b(p187), .O(EX465) );
and2 gate( .a(N165), .b(EX465), .O(EX466) );
and2 gate( .a(N451), .b(p188), .O(EX467) );
and2 gate( .a(N165), .b(EX467), .O(EX468) );
or2  gate( .a(EX462), .b(EX464), .O(EX469) );
or2  gate( .a(EX466), .b(EX469), .O(EX470) );
or2  gate( .a(EX468), .b(EX470), .O(N523) );
inv1 gate( .a(N451),.O(N451_NOT) );
inv1 gate( .a(N171),.O(N171_NOT));
and2 gate( .a(N451_NOT), .b(p189), .O(EX471) );
and2 gate( .a(N171_NOT), .b(EX471), .O(EX472) );
and2 gate( .a(N451), .b(p190), .O(EX473) );
and2 gate( .a(N171_NOT), .b(EX473), .O(EX474) );
and2 gate( .a(N451_NOT), .b(p191), .O(EX475) );
and2 gate( .a(N171), .b(EX475), .O(EX476) );
and2 gate( .a(N451), .b(p192), .O(EX477) );
and2 gate( .a(N171), .b(EX477), .O(EX478) );
or2  gate( .a(EX472), .b(EX474), .O(EX479) );
or2  gate( .a(EX476), .b(EX479), .O(EX480) );
or2  gate( .a(EX478), .b(EX480), .O(N524) );
inv1 gate( .a(N451),.O(N451_NOT) );
inv1 gate( .a(N177),.O(N177_NOT));
and2 gate( .a(N451_NOT), .b(p193), .O(EX481) );
and2 gate( .a(N177_NOT), .b(EX481), .O(EX482) );
and2 gate( .a(N451), .b(p194), .O(EX483) );
and2 gate( .a(N177_NOT), .b(EX483), .O(EX484) );
and2 gate( .a(N451_NOT), .b(p195), .O(EX485) );
and2 gate( .a(N177), .b(EX485), .O(EX486) );
and2 gate( .a(N451), .b(p196), .O(EX487) );
and2 gate( .a(N177), .b(EX487), .O(EX488) );
or2  gate( .a(EX482), .b(EX484), .O(EX489) );
or2  gate( .a(EX486), .b(EX489), .O(EX490) );
or2  gate( .a(EX488), .b(EX490), .O(N525) );
and2 gate172( .a(N451), .b(N183), .O(N526) );
nand2 gate173( .a(N451), .b(N189), .O(N527) );
inv1 gate( .a(N451),.O(N451_NOT) );
inv1 gate( .a(N195),.O(N195_NOT));
and2 gate( .a(N451_NOT), .b(p197), .O(EX491) );
and2 gate( .a(N195_NOT), .b(EX491), .O(EX492) );
and2 gate( .a(N451), .b(p198), .O(EX493) );
and2 gate( .a(N195_NOT), .b(EX493), .O(EX494) );
and2 gate( .a(N451_NOT), .b(p199), .O(EX495) );
and2 gate( .a(N195), .b(EX495), .O(EX496) );
and2 gate( .a(N451), .b(p200), .O(EX497) );
and2 gate( .a(N195), .b(EX497), .O(EX498) );
or2  gate( .a(EX492), .b(EX494), .O(EX499) );
or2  gate( .a(EX496), .b(EX499), .O(EX500) );
or2  gate( .a(EX498), .b(EX500), .O(N528) );
nand2 gate175( .a(N451), .b(N201), .O(N529) );
inv1 gate( .a(N498),.O(N498_NOT) );
inv1 gate( .a(N499),.O(N499_NOT));
and2 gate( .a(N498_NOT), .b(p201), .O(EX501) );
and2 gate( .a(N499_NOT), .b(EX501), .O(EX502) );
and2 gate( .a(N498), .b(p202), .O(EX503) );
and2 gate( .a(N499_NOT), .b(EX503), .O(EX504) );
and2 gate( .a(N498_NOT), .b(p203), .O(EX505) );
and2 gate( .a(N499), .b(EX505), .O(EX506) );
and2 gate( .a(N498), .b(p204), .O(EX507) );
and2 gate( .a(N499), .b(EX507), .O(EX508) );
or2  gate( .a(EX502), .b(EX504), .O(EX509) );
or2  gate( .a(EX506), .b(EX509), .O(EX510) );
or2  gate( .a(EX508), .b(EX510), .O(N530) );
nand2 gate177( .a(N500), .b(N501), .O(N533) );
nor2 gate178( .a(N309), .b(N502), .O(N536) );
nor2 gate179( .a(N316), .b(N504), .O(N537) );
inv1 gate( .a(N317),.O(N317_NOT) );
inv1 gate( .a(N506),.O(N506_NOT));
and2 gate( .a(N317_NOT), .b(p205), .O(EX511) );
and2 gate( .a(N506_NOT), .b(EX511), .O(EX512) );
and2 gate( .a(N317), .b(p206), .O(EX513) );
and2 gate( .a(N506_NOT), .b(EX513), .O(EX514) );
and2 gate( .a(N317_NOT), .b(p207), .O(EX515) );
and2 gate( .a(N506), .b(EX515), .O(EX516) );
and2 gate( .a(N317), .b(p208), .O(EX517) );
and2 gate( .a(N506), .b(EX517), .O(EX518) );
or2  gate( .a(EX512), .b(EX514), .O(EX519) );
or2  gate( .a(EX516), .b(EX519), .O(EX520) );
or2  gate( .a(EX518), .b(EX520), .O(N538) );
nor2 gate181( .a(N318), .b(N508), .O(N539) );
inv1 gate( .a(N510),.O(N510_NOT) );
inv1 gate( .a(N511),.O(N511_NOT));
and2 gate( .a(N510_NOT), .b(p209), .O(EX521) );
and2 gate( .a(N511_NOT), .b(EX521), .O(EX522) );
and2 gate( .a(N510), .b(p210), .O(EX523) );
and2 gate( .a(N511_NOT), .b(EX523), .O(EX524) );
and2 gate( .a(N510_NOT), .b(p211), .O(EX525) );
and2 gate( .a(N511), .b(EX525), .O(EX526) );
and2 gate( .a(N510), .b(p212), .O(EX527) );
and2 gate( .a(N511), .b(EX527), .O(EX528) );
or2  gate( .a(EX522), .b(EX524), .O(EX529) );
or2  gate( .a(EX526), .b(EX529), .O(EX530) );
or2  gate( .a(EX528), .b(EX530), .O(N540) );
nor2 gate183( .a(N512), .b(N513), .O(N541) );
inv1 gate( .a(N514),.O(N514_NOT) );
inv1 gate( .a(N515),.O(N515_NOT));
and2 gate( .a(N514_NOT), .b(p213), .O(EX531) );
and2 gate( .a(N515_NOT), .b(EX531), .O(EX532) );
and2 gate( .a(N514), .b(p214), .O(EX533) );
and2 gate( .a(N515_NOT), .b(EX533), .O(EX534) );
and2 gate( .a(N514_NOT), .b(p215), .O(EX535) );
and2 gate( .a(N515), .b(EX535), .O(EX536) );
and2 gate( .a(N514), .b(p216), .O(EX537) );
and2 gate( .a(N515), .b(EX537), .O(EX538) );
or2  gate( .a(EX532), .b(EX534), .O(EX539) );
or2  gate( .a(EX536), .b(EX539), .O(EX540) );
or2  gate( .a(EX538), .b(EX540), .O(N542) );
inv1 gate( .a(N516),.O(N516_NOT) );
inv1 gate( .a(N517),.O(N517_NOT));
and2 gate( .a(N516_NOT), .b(p217), .O(EX541) );
and2 gate( .a(N517_NOT), .b(EX541), .O(EX542) );
and2 gate( .a(N516), .b(p218), .O(EX543) );
and2 gate( .a(N517_NOT), .b(EX543), .O(EX544) );
and2 gate( .a(N516_NOT), .b(p219), .O(EX545) );
and2 gate( .a(N517), .b(EX545), .O(EX546) );
and2 gate( .a(N516), .b(p220), .O(EX547) );
and2 gate( .a(N517), .b(EX547), .O(EX548) );
or2  gate( .a(EX542), .b(EX544), .O(EX549) );
or2  gate( .a(EX546), .b(EX549), .O(EX550) );
or2  gate( .a(EX548), .b(EX550), .O(N543) );
inv1 gate( .a(N518),.O(N518_NOT) );
inv1 gate( .a(N519),.O(N519_NOT));
and2 gate( .a(N518_NOT), .b(p221), .O(EX551) );
and2 gate( .a(N519_NOT), .b(EX551), .O(EX552) );
and2 gate( .a(N518), .b(p222), .O(EX553) );
and2 gate( .a(N519_NOT), .b(EX553), .O(EX554) );
and2 gate( .a(N518_NOT), .b(p223), .O(EX555) );
and2 gate( .a(N519), .b(EX555), .O(EX556) );
and2 gate( .a(N518), .b(p224), .O(EX557) );
and2 gate( .a(N519), .b(EX557), .O(EX558) );
or2  gate( .a(EX552), .b(EX554), .O(EX559) );
or2  gate( .a(EX556), .b(EX559), .O(EX560) );
or2  gate( .a(EX558), .b(EX560), .O(N544) );
nand2 gate187( .a(N520), .b(N521), .O(N547) );
inv1 gate188( .a(N530), .O(N550) );
inv1 gate189( .a(N533), .O(N551) );
and2 gate190( .a(N530), .b(N533), .O(N552) );
nand2 gate191( .a(N536), .b(N503), .O(N553) );
nand2 gate192( .a(N537), .b(N505), .O(N557) );
nand2 gate193( .a(N538), .b(N507), .O(N561) );
nand2 gate194( .a(N539), .b(N509), .O(N565) );
inv1 gate( .a(N488),.O(N488_NOT) );
inv1 gate( .a(N540),.O(N540_NOT));
and2 gate( .a(N488_NOT), .b(p225), .O(EX561) );
and2 gate( .a(N540_NOT), .b(EX561), .O(EX562) );
and2 gate( .a(N488), .b(p226), .O(EX563) );
and2 gate( .a(N540_NOT), .b(EX563), .O(EX564) );
and2 gate( .a(N488_NOT), .b(p227), .O(EX565) );
and2 gate( .a(N540), .b(EX565), .O(EX566) );
and2 gate( .a(N488), .b(p228), .O(EX567) );
and2 gate( .a(N540), .b(EX567), .O(EX568) );
or2  gate( .a(EX562), .b(EX564), .O(EX569) );
or2  gate( .a(EX566), .b(EX569), .O(EX570) );
or2  gate( .a(EX568), .b(EX570), .O(N569) );
nand2 gate196( .a(N489), .b(N541), .O(N573) );
nand2 gate197( .a(N490), .b(N542), .O(N577) );
nand2 gate198( .a(N491), .b(N543), .O(N581) );
inv1 gate199( .a(N544), .O(N585) );
inv1 gate200( .a(N547), .O(N586) );
and2 gate201( .a(N544), .b(N547), .O(N587) );
inv1 gate( .a(N550),.O(N550_NOT) );
inv1 gate( .a(N551),.O(N551_NOT));
and2 gate( .a(N550_NOT), .b(p229), .O(EX571) );
and2 gate( .a(N551_NOT), .b(EX571), .O(EX572) );
and2 gate( .a(N550), .b(p230), .O(EX573) );
and2 gate( .a(N551_NOT), .b(EX573), .O(EX574) );
and2 gate( .a(N550_NOT), .b(p231), .O(EX575) );
and2 gate( .a(N551), .b(EX575), .O(EX576) );
and2 gate( .a(N550), .b(p232), .O(EX577) );
and2 gate( .a(N551), .b(EX577), .O(EX578) );
or2  gate( .a(EX572), .b(EX574), .O(EX579) );
or2  gate( .a(EX576), .b(EX579), .O(EX580) );
or2  gate( .a(EX578), .b(EX580), .O(N588) );
inv1 gate( .a(N585),.O(N585_NOT) );
inv1 gate( .a(N586),.O(N586_NOT));
and2 gate( .a(N585_NOT), .b(p233), .O(EX581) );
and2 gate( .a(N586_NOT), .b(EX581), .O(EX582) );
and2 gate( .a(N585), .b(p234), .O(EX583) );
and2 gate( .a(N586_NOT), .b(EX583), .O(EX584) );
and2 gate( .a(N585_NOT), .b(p235), .O(EX585) );
and2 gate( .a(N586), .b(EX585), .O(EX586) );
and2 gate( .a(N585), .b(p236), .O(EX587) );
and2 gate( .a(N586), .b(EX587), .O(EX588) );
or2  gate( .a(EX582), .b(EX584), .O(EX589) );
or2  gate( .a(EX586), .b(EX589), .O(EX590) );
or2  gate( .a(EX588), .b(EX590), .O(N589) );
inv1 gate( .a(N553),.O(N553_NOT) );
inv1 gate( .a(N159),.O(N159_NOT));
and2 gate( .a(N553_NOT), .b(p237), .O(EX591) );
and2 gate( .a(N159_NOT), .b(EX591), .O(EX592) );
and2 gate( .a(N553), .b(p238), .O(EX593) );
and2 gate( .a(N159_NOT), .b(EX593), .O(EX594) );
and2 gate( .a(N553_NOT), .b(p239), .O(EX595) );
and2 gate( .a(N159), .b(EX595), .O(EX596) );
and2 gate( .a(N553), .b(p240), .O(EX597) );
and2 gate( .a(N159), .b(EX597), .O(EX598) );
or2  gate( .a(EX592), .b(EX594), .O(EX599) );
or2  gate( .a(EX596), .b(EX599), .O(EX600) );
or2  gate( .a(EX598), .b(EX600), .O(N590) );
inv1 gate( .a(N553),.O(N553_NOT) );
inv1 gate( .a(N159),.O(N159_NOT));
and2 gate( .a(N553_NOT), .b(p241), .O(EX601) );
and2 gate( .a(N159_NOT), .b(EX601), .O(EX602) );
and2 gate( .a(N553), .b(p242), .O(EX603) );
and2 gate( .a(N159_NOT), .b(EX603), .O(EX604) );
and2 gate( .a(N553_NOT), .b(p243), .O(EX605) );
and2 gate( .a(N159), .b(EX605), .O(EX606) );
and2 gate( .a(N553), .b(p244), .O(EX607) );
and2 gate( .a(N159), .b(EX607), .O(EX608) );
or2  gate( .a(EX602), .b(EX604), .O(EX609) );
or2  gate( .a(EX606), .b(EX609), .O(EX610) );
or2  gate( .a(EX608), .b(EX610), .O(N593) );
and2 gate206( .a(N246), .b(N553), .O(N596) );
inv1 gate( .a(N557),.O(N557_NOT) );
inv1 gate( .a(N165),.O(N165_NOT));
and2 gate( .a(N557_NOT), .b(p245), .O(EX611) );
and2 gate( .a(N165_NOT), .b(EX611), .O(EX612) );
and2 gate( .a(N557), .b(p246), .O(EX613) );
and2 gate( .a(N165_NOT), .b(EX613), .O(EX614) );
and2 gate( .a(N557_NOT), .b(p247), .O(EX615) );
and2 gate( .a(N165), .b(EX615), .O(EX616) );
and2 gate( .a(N557), .b(p248), .O(EX617) );
and2 gate( .a(N165), .b(EX617), .O(EX618) );
or2  gate( .a(EX612), .b(EX614), .O(EX619) );
or2  gate( .a(EX616), .b(EX619), .O(EX620) );
or2  gate( .a(EX618), .b(EX620), .O(N597) );
or2 gate208( .a(N557), .b(N165), .O(N600) );
inv1 gate( .a(N246),.O(N246_NOT) );
inv1 gate( .a(N557),.O(N557_NOT));
and2 gate( .a(N246_NOT), .b(p249), .O(EX621) );
and2 gate( .a(N557_NOT), .b(EX621), .O(EX622) );
and2 gate( .a(N246), .b(p250), .O(EX623) );
and2 gate( .a(N557_NOT), .b(EX623), .O(EX624) );
and2 gate( .a(N246_NOT), .b(p251), .O(EX625) );
and2 gate( .a(N557), .b(EX625), .O(EX626) );
and2 gate( .a(N246), .b(p252), .O(EX627) );
and2 gate( .a(N557), .b(EX627), .O(EX628) );
or2  gate( .a(EX622), .b(EX624), .O(EX629) );
or2  gate( .a(EX626), .b(EX629), .O(EX630) );
or2  gate( .a(EX628), .b(EX630), .O(N605) );
inv1 gate( .a(N561),.O(N561_NOT) );
inv1 gate( .a(N171),.O(N171_NOT));
and2 gate( .a(N561_NOT), .b(p253), .O(EX631) );
and2 gate( .a(N171_NOT), .b(EX631), .O(EX632) );
and2 gate( .a(N561), .b(p254), .O(EX633) );
and2 gate( .a(N171_NOT), .b(EX633), .O(EX634) );
and2 gate( .a(N561_NOT), .b(p255), .O(EX635) );
and2 gate( .a(N171), .b(EX635), .O(EX636) );
and2 gate( .a(N561), .b(p256), .O(EX637) );
and2 gate( .a(N171), .b(EX637), .O(EX638) );
or2  gate( .a(EX632), .b(EX634), .O(EX639) );
or2  gate( .a(EX636), .b(EX639), .O(EX640) );
or2  gate( .a(EX638), .b(EX640), .O(N606) );
or2 gate211( .a(N561), .b(N171), .O(N609) );
and2 gate212( .a(N246), .b(N561), .O(N615) );
nand2 gate213( .a(N565), .b(N177), .O(N616) );
inv1 gate( .a(N565),.O(N565_NOT) );
inv1 gate( .a(N177),.O(N177_NOT));
and2 gate( .a(N565_NOT), .b(p257), .O(EX641) );
and2 gate( .a(N177_NOT), .b(EX641), .O(EX642) );
and2 gate( .a(N565), .b(p258), .O(EX643) );
and2 gate( .a(N177_NOT), .b(EX643), .O(EX644) );
and2 gate( .a(N565_NOT), .b(p259), .O(EX645) );
and2 gate( .a(N177), .b(EX645), .O(EX646) );
and2 gate( .a(N565), .b(p260), .O(EX647) );
and2 gate( .a(N177), .b(EX647), .O(EX648) );
or2  gate( .a(EX642), .b(EX644), .O(EX649) );
or2  gate( .a(EX646), .b(EX649), .O(EX650) );
or2  gate( .a(EX648), .b(EX650), .O(N619) );
and2 gate215( .a(N246), .b(N565), .O(N624) );
inv1 gate( .a(N569),.O(N569_NOT) );
inv1 gate( .a(N183),.O(N183_NOT));
and2 gate( .a(N569_NOT), .b(p261), .O(EX651) );
and2 gate( .a(N183_NOT), .b(EX651), .O(EX652) );
and2 gate( .a(N569), .b(p262), .O(EX653) );
and2 gate( .a(N183_NOT), .b(EX653), .O(EX654) );
and2 gate( .a(N569_NOT), .b(p263), .O(EX655) );
and2 gate( .a(N183), .b(EX655), .O(EX656) );
and2 gate( .a(N569), .b(p264), .O(EX657) );
and2 gate( .a(N183), .b(EX657), .O(EX658) );
or2  gate( .a(EX652), .b(EX654), .O(EX659) );
or2  gate( .a(EX656), .b(EX659), .O(EX660) );
or2  gate( .a(EX658), .b(EX660), .O(N625) );
inv1 gate( .a(N569),.O(N569_NOT) );
inv1 gate( .a(N183),.O(N183_NOT));
and2 gate( .a(N569_NOT), .b(p265), .O(EX661) );
and2 gate( .a(N183_NOT), .b(EX661), .O(EX662) );
and2 gate( .a(N569), .b(p266), .O(EX663) );
and2 gate( .a(N183_NOT), .b(EX663), .O(EX664) );
and2 gate( .a(N569_NOT), .b(p267), .O(EX665) );
and2 gate( .a(N183), .b(EX665), .O(EX666) );
and2 gate( .a(N569), .b(p268), .O(EX667) );
and2 gate( .a(N183), .b(EX667), .O(EX668) );
or2  gate( .a(EX662), .b(EX664), .O(EX669) );
or2  gate( .a(EX666), .b(EX669), .O(EX670) );
or2  gate( .a(EX668), .b(EX670), .O(N628) );
inv1 gate( .a(N246),.O(N246_NOT) );
inv1 gate( .a(N569),.O(N569_NOT));
and2 gate( .a(N246_NOT), .b(p269), .O(EX671) );
and2 gate( .a(N569_NOT), .b(EX671), .O(EX672) );
and2 gate( .a(N246), .b(p270), .O(EX673) );
and2 gate( .a(N569_NOT), .b(EX673), .O(EX674) );
and2 gate( .a(N246_NOT), .b(p271), .O(EX675) );
and2 gate( .a(N569), .b(EX675), .O(EX676) );
and2 gate( .a(N246), .b(p272), .O(EX677) );
and2 gate( .a(N569), .b(EX677), .O(EX678) );
or2  gate( .a(EX672), .b(EX674), .O(EX679) );
or2  gate( .a(EX676), .b(EX679), .O(EX680) );
or2  gate( .a(EX678), .b(EX680), .O(N631) );
nand2 gate219( .a(N573), .b(N189), .O(N632) );
inv1 gate( .a(N573),.O(N573_NOT) );
inv1 gate( .a(N189),.O(N189_NOT));
and2 gate( .a(N573_NOT), .b(p273), .O(EX681) );
and2 gate( .a(N189_NOT), .b(EX681), .O(EX682) );
and2 gate( .a(N573), .b(p274), .O(EX683) );
and2 gate( .a(N189_NOT), .b(EX683), .O(EX684) );
and2 gate( .a(N573_NOT), .b(p275), .O(EX685) );
and2 gate( .a(N189), .b(EX685), .O(EX686) );
and2 gate( .a(N573), .b(p276), .O(EX687) );
and2 gate( .a(N189), .b(EX687), .O(EX688) );
or2  gate( .a(EX682), .b(EX684), .O(EX689) );
or2  gate( .a(EX686), .b(EX689), .O(EX690) );
or2  gate( .a(EX688), .b(EX690), .O(N635) );
and2 gate221( .a(N246), .b(N573), .O(N640) );
nand2 gate222( .a(N577), .b(N195), .O(N641) );
or2 gate223( .a(N577), .b(N195), .O(N644) );
and2 gate224( .a(N246), .b(N577), .O(N650) );
nand2 gate225( .a(N581), .b(N201), .O(N651) );
inv1 gate( .a(N581),.O(N581_NOT) );
inv1 gate( .a(N201),.O(N201_NOT));
and2 gate( .a(N581_NOT), .b(p277), .O(EX691) );
and2 gate( .a(N201_NOT), .b(EX691), .O(EX692) );
and2 gate( .a(N581), .b(p278), .O(EX693) );
and2 gate( .a(N201_NOT), .b(EX693), .O(EX694) );
and2 gate( .a(N581_NOT), .b(p279), .O(EX695) );
and2 gate( .a(N201), .b(EX695), .O(EX696) );
and2 gate( .a(N581), .b(p280), .O(EX697) );
and2 gate( .a(N201), .b(EX697), .O(EX698) );
or2  gate( .a(EX692), .b(EX694), .O(EX699) );
or2  gate( .a(EX696), .b(EX699), .O(EX700) );
or2  gate( .a(EX698), .b(EX700), .O(N654) );
inv1 gate( .a(N246),.O(N246_NOT) );
inv1 gate( .a(N581),.O(N581_NOT));
and2 gate( .a(N246_NOT), .b(p281), .O(EX701) );
and2 gate( .a(N581_NOT), .b(EX701), .O(EX702) );
and2 gate( .a(N246), .b(p282), .O(EX703) );
and2 gate( .a(N581_NOT), .b(EX703), .O(EX704) );
and2 gate( .a(N246_NOT), .b(p283), .O(EX705) );
and2 gate( .a(N581), .b(EX705), .O(EX706) );
and2 gate( .a(N246), .b(p284), .O(EX707) );
and2 gate( .a(N581), .b(EX707), .O(EX708) );
or2  gate( .a(EX702), .b(EX704), .O(EX709) );
or2  gate( .a(EX706), .b(EX709), .O(EX710) );
or2  gate( .a(EX708), .b(EX710), .O(N659) );
nor2 gate228( .a(N552), .b(N588), .O(N660) );
inv1 gate( .a(N587),.O(N587_NOT) );
inv1 gate( .a(N589),.O(N589_NOT));
and2 gate( .a(N587_NOT), .b(p285), .O(EX711) );
and2 gate( .a(N589_NOT), .b(EX711), .O(EX712) );
and2 gate( .a(N587), .b(p286), .O(EX713) );
and2 gate( .a(N589_NOT), .b(EX713), .O(EX714) );
and2 gate( .a(N587_NOT), .b(p287), .O(EX715) );
and2 gate( .a(N589), .b(EX715), .O(EX716) );
and2 gate( .a(N587), .b(p288), .O(EX717) );
and2 gate( .a(N589), .b(EX717), .O(EX718) );
or2  gate( .a(EX712), .b(EX714), .O(EX719) );
or2  gate( .a(EX716), .b(EX719), .O(EX720) );
or2  gate( .a(EX718), .b(EX720), .O(N661) );
inv1 gate230( .a(N590), .O(N662) );
inv1 gate( .a(N593),.O(N593_NOT) );
inv1 gate( .a(N590),.O(N590_NOT));
and2 gate( .a(N593_NOT), .b(p289), .O(EX721) );
and2 gate( .a(N590_NOT), .b(EX721), .O(EX722) );
and2 gate( .a(N593), .b(p290), .O(EX723) );
and2 gate( .a(N590_NOT), .b(EX723), .O(EX724) );
and2 gate( .a(N593_NOT), .b(p291), .O(EX725) );
and2 gate( .a(N590), .b(EX725), .O(EX726) );
and2 gate( .a(N593), .b(p292), .O(EX727) );
and2 gate( .a(N590), .b(EX727), .O(EX728) );
or2  gate( .a(EX722), .b(EX724), .O(EX729) );
or2  gate( .a(EX726), .b(EX729), .O(EX730) );
or2  gate( .a(EX728), .b(EX730), .O(N665) );
inv1 gate( .a(N596),.O(N596_NOT) );
inv1 gate( .a(N522),.O(N522_NOT));
and2 gate( .a(N596_NOT), .b(p293), .O(EX731) );
and2 gate( .a(N522_NOT), .b(EX731), .O(EX732) );
and2 gate( .a(N596), .b(p294), .O(EX733) );
and2 gate( .a(N522_NOT), .b(EX733), .O(EX734) );
and2 gate( .a(N596_NOT), .b(p295), .O(EX735) );
and2 gate( .a(N522), .b(EX735), .O(EX736) );
and2 gate( .a(N596), .b(p296), .O(EX737) );
and2 gate( .a(N522), .b(EX737), .O(EX738) );
or2  gate( .a(EX732), .b(EX734), .O(EX739) );
or2  gate( .a(EX736), .b(EX739), .O(EX740) );
or2  gate( .a(EX738), .b(EX740), .O(N669) );
inv1 gate233( .a(N597), .O(N670) );
and2 gate234( .a(N600), .b(N597), .O(N673) );
nor2 gate235( .a(N605), .b(N523), .O(N677) );
inv1 gate236( .a(N606), .O(N678) );
inv1 gate( .a(N609),.O(N609_NOT) );
inv1 gate( .a(N606),.O(N606_NOT));
and2 gate( .a(N609_NOT), .b(p297), .O(EX741) );
and2 gate( .a(N606_NOT), .b(EX741), .O(EX742) );
and2 gate( .a(N609), .b(p298), .O(EX743) );
and2 gate( .a(N606_NOT), .b(EX743), .O(EX744) );
and2 gate( .a(N609_NOT), .b(p299), .O(EX745) );
and2 gate( .a(N606), .b(EX745), .O(EX746) );
and2 gate( .a(N609), .b(p300), .O(EX747) );
and2 gate( .a(N606), .b(EX747), .O(EX748) );
or2  gate( .a(EX742), .b(EX744), .O(EX749) );
or2  gate( .a(EX746), .b(EX749), .O(EX750) );
or2  gate( .a(EX748), .b(EX750), .O(N682) );
nor2 gate238( .a(N615), .b(N524), .O(N686) );
inv1 gate239( .a(N616), .O(N687) );
and2 gate240( .a(N619), .b(N616), .O(N692) );
nor2 gate241( .a(N624), .b(N525), .O(N696) );
inv1 gate242( .a(N625), .O(N697) );
and2 gate243( .a(N628), .b(N625), .O(N700) );
inv1 gate( .a(N631),.O(N631_NOT) );
inv1 gate( .a(N526),.O(N526_NOT));
and2 gate( .a(N631_NOT), .b(p301), .O(EX751) );
and2 gate( .a(N526_NOT), .b(EX751), .O(EX752) );
and2 gate( .a(N631), .b(p302), .O(EX753) );
and2 gate( .a(N526_NOT), .b(EX753), .O(EX754) );
and2 gate( .a(N631_NOT), .b(p303), .O(EX755) );
and2 gate( .a(N526), .b(EX755), .O(EX756) );
and2 gate( .a(N631), .b(p304), .O(EX757) );
and2 gate( .a(N526), .b(EX757), .O(EX758) );
or2  gate( .a(EX752), .b(EX754), .O(EX759) );
or2  gate( .a(EX756), .b(EX759), .O(EX760) );
or2  gate( .a(EX758), .b(EX760), .O(N704) );
inv1 gate245( .a(N632), .O(N705) );
inv1 gate( .a(N635),.O(N635_NOT) );
inv1 gate( .a(N632),.O(N632_NOT));
and2 gate( .a(N635_NOT), .b(p305), .O(EX761) );
and2 gate( .a(N632_NOT), .b(EX761), .O(EX762) );
and2 gate( .a(N635), .b(p306), .O(EX763) );
and2 gate( .a(N632_NOT), .b(EX763), .O(EX764) );
and2 gate( .a(N635_NOT), .b(p307), .O(EX765) );
and2 gate( .a(N632), .b(EX765), .O(EX766) );
and2 gate( .a(N635), .b(p308), .O(EX767) );
and2 gate( .a(N632), .b(EX767), .O(EX768) );
or2  gate( .a(EX762), .b(EX764), .O(EX769) );
or2  gate( .a(EX766), .b(EX769), .O(EX770) );
or2  gate( .a(EX768), .b(EX770), .O(N708) );
nor2 gate247( .a(N337), .b(N640), .O(N712) );
inv1 gate248( .a(N641), .O(N713) );
and2 gate249( .a(N644), .b(N641), .O(N717) );
nor2 gate250( .a(N339), .b(N650), .O(N721) );
inv1 gate251( .a(N651), .O(N722) );
inv1 gate( .a(N654),.O(N654_NOT) );
inv1 gate( .a(N651),.O(N651_NOT));
and2 gate( .a(N654_NOT), .b(p309), .O(EX771) );
and2 gate( .a(N651_NOT), .b(EX771), .O(EX772) );
and2 gate( .a(N654), .b(p310), .O(EX773) );
and2 gate( .a(N651_NOT), .b(EX773), .O(EX774) );
and2 gate( .a(N654_NOT), .b(p311), .O(EX775) );
and2 gate( .a(N651), .b(EX775), .O(EX776) );
and2 gate( .a(N654), .b(p312), .O(EX777) );
and2 gate( .a(N651), .b(EX777), .O(EX778) );
or2  gate( .a(EX772), .b(EX774), .O(EX779) );
or2  gate( .a(EX776), .b(EX779), .O(EX780) );
or2  gate( .a(EX778), .b(EX780), .O(N727) );
nor2 gate253( .a(N341), .b(N659), .O(N731) );
nand2 gate254( .a(N654), .b(N261), .O(N732) );
nand3 gate255( .a(N644), .b(N654), .c(N261), .O(N733) );
nand4 gate256( .a(N635), .b(N644), .c(N654), .d(N261), .O(N734) );
inv1 gate257( .a(N662), .O(N735) );
inv1 gate( .a(N228),.O(N228_NOT) );
inv1 gate( .a(N665),.O(N665_NOT));
and2 gate( .a(N228_NOT), .b(p313), .O(EX781) );
and2 gate( .a(N665_NOT), .b(EX781), .O(EX782) );
and2 gate( .a(N228), .b(p314), .O(EX783) );
and2 gate( .a(N665_NOT), .b(EX783), .O(EX784) );
and2 gate( .a(N228_NOT), .b(p315), .O(EX785) );
and2 gate( .a(N665), .b(EX785), .O(EX786) );
and2 gate( .a(N228), .b(p316), .O(EX787) );
and2 gate( .a(N665), .b(EX787), .O(EX788) );
or2  gate( .a(EX782), .b(EX784), .O(EX789) );
or2  gate( .a(EX786), .b(EX789), .O(EX790) );
or2  gate( .a(EX788), .b(EX790), .O(N736) );
inv1 gate( .a(N237),.O(N237_NOT) );
inv1 gate( .a(N662),.O(N662_NOT));
and2 gate( .a(N237_NOT), .b(p317), .O(EX791) );
and2 gate( .a(N662_NOT), .b(EX791), .O(EX792) );
and2 gate( .a(N237), .b(p318), .O(EX793) );
and2 gate( .a(N662_NOT), .b(EX793), .O(EX794) );
and2 gate( .a(N237_NOT), .b(p319), .O(EX795) );
and2 gate( .a(N662), .b(EX795), .O(EX796) );
and2 gate( .a(N237), .b(p320), .O(EX797) );
and2 gate( .a(N662), .b(EX797), .O(EX798) );
or2  gate( .a(EX792), .b(EX794), .O(EX799) );
or2  gate( .a(EX796), .b(EX799), .O(EX800) );
or2  gate( .a(EX798), .b(EX800), .O(N737) );
inv1 gate260( .a(N670), .O(N738) );
and2 gate261( .a(N228), .b(N673), .O(N739) );
and2 gate262( .a(N237), .b(N670), .O(N740) );
inv1 gate263( .a(N678), .O(N741) );
inv1 gate( .a(N228),.O(N228_NOT) );
inv1 gate( .a(N682),.O(N682_NOT));
and2 gate( .a(N228_NOT), .b(p321), .O(EX801) );
and2 gate( .a(N682_NOT), .b(EX801), .O(EX802) );
and2 gate( .a(N228), .b(p322), .O(EX803) );
and2 gate( .a(N682_NOT), .b(EX803), .O(EX804) );
and2 gate( .a(N228_NOT), .b(p323), .O(EX805) );
and2 gate( .a(N682), .b(EX805), .O(EX806) );
and2 gate( .a(N228), .b(p324), .O(EX807) );
and2 gate( .a(N682), .b(EX807), .O(EX808) );
or2  gate( .a(EX802), .b(EX804), .O(EX809) );
or2  gate( .a(EX806), .b(EX809), .O(EX810) );
or2  gate( .a(EX808), .b(EX810), .O(N742) );
inv1 gate( .a(N237),.O(N237_NOT) );
inv1 gate( .a(N678),.O(N678_NOT));
and2 gate( .a(N237_NOT), .b(p325), .O(EX811) );
and2 gate( .a(N678_NOT), .b(EX811), .O(EX812) );
and2 gate( .a(N237), .b(p326), .O(EX813) );
and2 gate( .a(N678_NOT), .b(EX813), .O(EX814) );
and2 gate( .a(N237_NOT), .b(p327), .O(EX815) );
and2 gate( .a(N678), .b(EX815), .O(EX816) );
and2 gate( .a(N237), .b(p328), .O(EX817) );
and2 gate( .a(N678), .b(EX817), .O(EX818) );
or2  gate( .a(EX812), .b(EX814), .O(EX819) );
or2  gate( .a(EX816), .b(EX819), .O(EX820) );
or2  gate( .a(EX818), .b(EX820), .O(N743) );
inv1 gate266( .a(N687), .O(N744) );
and2 gate267( .a(N228), .b(N692), .O(N745) );
inv1 gate( .a(N237),.O(N237_NOT) );
inv1 gate( .a(N687),.O(N687_NOT));
and2 gate( .a(N237_NOT), .b(p329), .O(EX821) );
and2 gate( .a(N687_NOT), .b(EX821), .O(EX822) );
and2 gate( .a(N237), .b(p330), .O(EX823) );
and2 gate( .a(N687_NOT), .b(EX823), .O(EX824) );
and2 gate( .a(N237_NOT), .b(p331), .O(EX825) );
and2 gate( .a(N687), .b(EX825), .O(EX826) );
and2 gate( .a(N237), .b(p332), .O(EX827) );
and2 gate( .a(N687), .b(EX827), .O(EX828) );
or2  gate( .a(EX822), .b(EX824), .O(EX829) );
or2  gate( .a(EX826), .b(EX829), .O(EX830) );
or2  gate( .a(EX828), .b(EX830), .O(N746) );
inv1 gate269( .a(N697), .O(N747) );
inv1 gate( .a(N228),.O(N228_NOT) );
inv1 gate( .a(N700),.O(N700_NOT));
and2 gate( .a(N228_NOT), .b(p333), .O(EX831) );
and2 gate( .a(N700_NOT), .b(EX831), .O(EX832) );
and2 gate( .a(N228), .b(p334), .O(EX833) );
and2 gate( .a(N700_NOT), .b(EX833), .O(EX834) );
and2 gate( .a(N228_NOT), .b(p335), .O(EX835) );
and2 gate( .a(N700), .b(EX835), .O(EX836) );
and2 gate( .a(N228), .b(p336), .O(EX837) );
and2 gate( .a(N700), .b(EX837), .O(EX838) );
or2  gate( .a(EX832), .b(EX834), .O(EX839) );
or2  gate( .a(EX836), .b(EX839), .O(EX840) );
or2  gate( .a(EX838), .b(EX840), .O(N748) );
and2 gate271( .a(N237), .b(N697), .O(N749) );
inv1 gate272( .a(N705), .O(N750) );
inv1 gate( .a(N228),.O(N228_NOT) );
inv1 gate( .a(N708),.O(N708_NOT));
and2 gate( .a(N228_NOT), .b(p337), .O(EX841) );
and2 gate( .a(N708_NOT), .b(EX841), .O(EX842) );
and2 gate( .a(N228), .b(p338), .O(EX843) );
and2 gate( .a(N708_NOT), .b(EX843), .O(EX844) );
and2 gate( .a(N228_NOT), .b(p339), .O(EX845) );
and2 gate( .a(N708), .b(EX845), .O(EX846) );
and2 gate( .a(N228), .b(p340), .O(EX847) );
and2 gate( .a(N708), .b(EX847), .O(EX848) );
or2  gate( .a(EX842), .b(EX844), .O(EX849) );
or2  gate( .a(EX846), .b(EX849), .O(EX850) );
or2  gate( .a(EX848), .b(EX850), .O(N751) );
and2 gate274( .a(N237), .b(N705), .O(N752) );
inv1 gate275( .a(N713), .O(N753) );
and2 gate276( .a(N228), .b(N717), .O(N754) );
inv1 gate( .a(N237),.O(N237_NOT) );
inv1 gate( .a(N713),.O(N713_NOT));
and2 gate( .a(N237_NOT), .b(p341), .O(EX851) );
and2 gate( .a(N713_NOT), .b(EX851), .O(EX852) );
and2 gate( .a(N237), .b(p342), .O(EX853) );
and2 gate( .a(N713_NOT), .b(EX853), .O(EX854) );
and2 gate( .a(N237_NOT), .b(p343), .O(EX855) );
and2 gate( .a(N713), .b(EX855), .O(EX856) );
and2 gate( .a(N237), .b(p344), .O(EX857) );
and2 gate( .a(N713), .b(EX857), .O(EX858) );
or2  gate( .a(EX852), .b(EX854), .O(EX859) );
or2  gate( .a(EX856), .b(EX859), .O(EX860) );
or2  gate( .a(EX858), .b(EX860), .O(N755) );
inv1 gate278( .a(N722), .O(N756) );
nor2 gate279( .a(N727), .b(N261), .O(N757) );
and2 gate280( .a(N727), .b(N261), .O(N758) );
inv1 gate( .a(N228),.O(N228_NOT) );
inv1 gate( .a(N727),.O(N727_NOT));
and2 gate( .a(N228_NOT), .b(p345), .O(EX861) );
and2 gate( .a(N727_NOT), .b(EX861), .O(EX862) );
and2 gate( .a(N228), .b(p346), .O(EX863) );
and2 gate( .a(N727_NOT), .b(EX863), .O(EX864) );
and2 gate( .a(N228_NOT), .b(p347), .O(EX865) );
and2 gate( .a(N727), .b(EX865), .O(EX866) );
and2 gate( .a(N228), .b(p348), .O(EX867) );
and2 gate( .a(N727), .b(EX867), .O(EX868) );
or2  gate( .a(EX862), .b(EX864), .O(EX869) );
or2  gate( .a(EX866), .b(EX869), .O(EX870) );
or2  gate( .a(EX868), .b(EX870), .O(N759) );
and2 gate282( .a(N237), .b(N722), .O(N760) );
nand2 gate283( .a(N644), .b(N722), .O(N761) );
nand2 gate284( .a(N635), .b(N713), .O(N762) );
nand3 gate285( .a(N635), .b(N644), .c(N722), .O(N763) );
nand2 gate286( .a(N609), .b(N687), .O(N764) );
inv1 gate( .a(N600),.O(N600_NOT) );
inv1 gate( .a(N678),.O(N678_NOT));
and2 gate( .a(N600_NOT), .b(p349), .O(EX871) );
and2 gate( .a(N678_NOT), .b(EX871), .O(EX872) );
and2 gate( .a(N600), .b(p350), .O(EX873) );
and2 gate( .a(N678_NOT), .b(EX873), .O(EX874) );
and2 gate( .a(N600_NOT), .b(p351), .O(EX875) );
and2 gate( .a(N678), .b(EX875), .O(EX876) );
and2 gate( .a(N600), .b(p352), .O(EX877) );
and2 gate( .a(N678), .b(EX877), .O(EX878) );
or2  gate( .a(EX872), .b(EX874), .O(EX879) );
or2  gate( .a(EX876), .b(EX879), .O(EX880) );
or2  gate( .a(EX878), .b(EX880), .O(N765) );
nand3 gate288( .a(N600), .b(N609), .c(N687), .O(N766) );
buf1 gate289( .a(N660), .O(N767) );
buf1 gate290( .a(N661), .O(N768) );
inv1 gate( .a(N736),.O(N736_NOT) );
inv1 gate( .a(N737),.O(N737_NOT));
and2 gate( .a(N736_NOT), .b(p353), .O(EX881) );
and2 gate( .a(N737_NOT), .b(EX881), .O(EX882) );
and2 gate( .a(N736), .b(p354), .O(EX883) );
and2 gate( .a(N737_NOT), .b(EX883), .O(EX884) );
and2 gate( .a(N736_NOT), .b(p355), .O(EX885) );
and2 gate( .a(N737), .b(EX885), .O(EX886) );
and2 gate( .a(N736), .b(p356), .O(EX887) );
and2 gate( .a(N737), .b(EX887), .O(EX888) );
or2  gate( .a(EX882), .b(EX884), .O(EX889) );
or2  gate( .a(EX886), .b(EX889), .O(EX890) );
or2  gate( .a(EX888), .b(EX890), .O(N769) );
nor2 gate292( .a(N739), .b(N740), .O(N770) );
nor2 gate293( .a(N742), .b(N743), .O(N771) );
nor2 gate294( .a(N745), .b(N746), .O(N772) );
nand4 gate295( .a(N750), .b(N762), .c(N763), .d(N734), .O(N773) );
inv1 gate( .a(N748),.O(N748_NOT) );
inv1 gate( .a(N749),.O(N749_NOT));
and2 gate( .a(N748_NOT), .b(p357), .O(EX891) );
and2 gate( .a(N749_NOT), .b(EX891), .O(EX892) );
and2 gate( .a(N748), .b(p358), .O(EX893) );
and2 gate( .a(N749_NOT), .b(EX893), .O(EX894) );
and2 gate( .a(N748_NOT), .b(p359), .O(EX895) );
and2 gate( .a(N749), .b(EX895), .O(EX896) );
and2 gate( .a(N748), .b(p360), .O(EX897) );
and2 gate( .a(N749), .b(EX897), .O(EX898) );
or2  gate( .a(EX892), .b(EX894), .O(EX899) );
or2  gate( .a(EX896), .b(EX899), .O(EX900) );
or2  gate( .a(EX898), .b(EX900), .O(N777) );
nand3 gate297( .a(N753), .b(N761), .c(N733), .O(N778) );
inv1 gate( .a(N751),.O(N751_NOT) );
inv1 gate( .a(N752),.O(N752_NOT));
and2 gate( .a(N751_NOT), .b(p361), .O(EX901) );
and2 gate( .a(N752_NOT), .b(EX901), .O(EX902) );
and2 gate( .a(N751), .b(p362), .O(EX903) );
and2 gate( .a(N752_NOT), .b(EX903), .O(EX904) );
and2 gate( .a(N751_NOT), .b(p363), .O(EX905) );
and2 gate( .a(N752), .b(EX905), .O(EX906) );
and2 gate( .a(N751), .b(p364), .O(EX907) );
and2 gate( .a(N752), .b(EX907), .O(EX908) );
or2  gate( .a(EX902), .b(EX904), .O(EX909) );
or2  gate( .a(EX906), .b(EX909), .O(EX910) );
or2  gate( .a(EX908), .b(EX910), .O(N781) );
inv1 gate( .a(N756),.O(N756_NOT) );
inv1 gate( .a(N732),.O(N732_NOT));
and2 gate( .a(N756_NOT), .b(p365), .O(EX911) );
and2 gate( .a(N732_NOT), .b(EX911), .O(EX912) );
and2 gate( .a(N756), .b(p366), .O(EX913) );
and2 gate( .a(N732_NOT), .b(EX913), .O(EX914) );
and2 gate( .a(N756_NOT), .b(p367), .O(EX915) );
and2 gate( .a(N732), .b(EX915), .O(EX916) );
and2 gate( .a(N756), .b(p368), .O(EX917) );
and2 gate( .a(N732), .b(EX917), .O(EX918) );
or2  gate( .a(EX912), .b(EX914), .O(EX919) );
or2  gate( .a(EX916), .b(EX919), .O(EX920) );
or2  gate( .a(EX918), .b(EX920), .O(N782) );
inv1 gate( .a(N754),.O(N754_NOT) );
inv1 gate( .a(N755),.O(N755_NOT));
and2 gate( .a(N754_NOT), .b(p369), .O(EX921) );
and2 gate( .a(N755_NOT), .b(EX921), .O(EX922) );
and2 gate( .a(N754), .b(p370), .O(EX923) );
and2 gate( .a(N755_NOT), .b(EX923), .O(EX924) );
and2 gate( .a(N754_NOT), .b(p371), .O(EX925) );
and2 gate( .a(N755), .b(EX925), .O(EX926) );
and2 gate( .a(N754), .b(p372), .O(EX927) );
and2 gate( .a(N755), .b(EX927), .O(EX928) );
or2  gate( .a(EX922), .b(EX924), .O(EX929) );
or2  gate( .a(EX926), .b(EX929), .O(EX930) );
or2  gate( .a(EX928), .b(EX930), .O(N785) );
nor2 gate301( .a(N757), .b(N758), .O(N786) );
nor2 gate302( .a(N759), .b(N760), .O(N787) );
inv1 gate( .a(N700),.O(N700_NOT) );
inv1 gate( .a(N773),.O(N773_NOT));
and2 gate( .a(N700_NOT), .b(p373), .O(EX931) );
and2 gate( .a(N773_NOT), .b(EX931), .O(EX932) );
and2 gate( .a(N700), .b(p374), .O(EX933) );
and2 gate( .a(N773_NOT), .b(EX933), .O(EX934) );
and2 gate( .a(N700_NOT), .b(p375), .O(EX935) );
and2 gate( .a(N773), .b(EX935), .O(EX936) );
and2 gate( .a(N700), .b(p376), .O(EX937) );
and2 gate( .a(N773), .b(EX937), .O(EX938) );
or2  gate( .a(EX932), .b(EX934), .O(EX939) );
or2  gate( .a(EX936), .b(EX939), .O(EX940) );
or2  gate( .a(EX938), .b(EX940), .O(N788) );
inv1 gate( .a(N700),.O(N700_NOT) );
inv1 gate( .a(N773),.O(N773_NOT));
and2 gate( .a(N700_NOT), .b(p377), .O(EX941) );
and2 gate( .a(N773_NOT), .b(EX941), .O(EX942) );
and2 gate( .a(N700), .b(p378), .O(EX943) );
and2 gate( .a(N773_NOT), .b(EX943), .O(EX944) );
and2 gate( .a(N700_NOT), .b(p379), .O(EX945) );
and2 gate( .a(N773), .b(EX945), .O(EX946) );
and2 gate( .a(N700), .b(p380), .O(EX947) );
and2 gate( .a(N773), .b(EX947), .O(EX948) );
or2  gate( .a(EX942), .b(EX944), .O(EX949) );
or2  gate( .a(EX946), .b(EX949), .O(EX950) );
or2  gate( .a(EX948), .b(EX950), .O(N789) );
inv1 gate( .a(N708),.O(N708_NOT) );
inv1 gate( .a(N778),.O(N778_NOT));
and2 gate( .a(N708_NOT), .b(p381), .O(EX951) );
and2 gate( .a(N778_NOT), .b(EX951), .O(EX952) );
and2 gate( .a(N708), .b(p382), .O(EX953) );
and2 gate( .a(N778_NOT), .b(EX953), .O(EX954) );
and2 gate( .a(N708_NOT), .b(p383), .O(EX955) );
and2 gate( .a(N778), .b(EX955), .O(EX956) );
and2 gate( .a(N708), .b(p384), .O(EX957) );
and2 gate( .a(N778), .b(EX957), .O(EX958) );
or2  gate( .a(EX952), .b(EX954), .O(EX959) );
or2  gate( .a(EX956), .b(EX959), .O(EX960) );
or2  gate( .a(EX958), .b(EX960), .O(N790) );
and2 gate306( .a(N708), .b(N778), .O(N791) );
nor2 gate307( .a(N717), .b(N782), .O(N792) );
and2 gate308( .a(N717), .b(N782), .O(N793) );
and2 gate309( .a(N219), .b(N786), .O(N794) );
inv1 gate( .a(N628),.O(N628_NOT) );
inv1 gate( .a(N773),.O(N773_NOT));
and2 gate( .a(N628_NOT), .b(p385), .O(EX961) );
and2 gate( .a(N773_NOT), .b(EX961), .O(EX962) );
and2 gate( .a(N628), .b(p386), .O(EX963) );
and2 gate( .a(N773_NOT), .b(EX963), .O(EX964) );
and2 gate( .a(N628_NOT), .b(p387), .O(EX965) );
and2 gate( .a(N773), .b(EX965), .O(EX966) );
and2 gate( .a(N628), .b(p388), .O(EX967) );
and2 gate( .a(N773), .b(EX967), .O(EX968) );
or2  gate( .a(EX962), .b(EX964), .O(EX969) );
or2  gate( .a(EX966), .b(EX969), .O(EX970) );
or2  gate( .a(EX968), .b(EX970), .O(N795) );
inv1 gate( .a(N795),.O(N795_NOT) );
inv1 gate( .a(N747),.O(N747_NOT));
and2 gate( .a(N795_NOT), .b(p389), .O(EX971) );
and2 gate( .a(N747_NOT), .b(EX971), .O(EX972) );
and2 gate( .a(N795), .b(p390), .O(EX973) );
and2 gate( .a(N747_NOT), .b(EX973), .O(EX974) );
and2 gate( .a(N795_NOT), .b(p391), .O(EX975) );
and2 gate( .a(N747), .b(EX975), .O(EX976) );
and2 gate( .a(N795), .b(p392), .O(EX977) );
and2 gate( .a(N747), .b(EX977), .O(EX978) );
or2  gate( .a(EX972), .b(EX974), .O(EX979) );
or2  gate( .a(EX976), .b(EX979), .O(EX980) );
or2  gate( .a(EX978), .b(EX980), .O(N796) );
inv1 gate( .a(N788),.O(N788_NOT) );
inv1 gate( .a(N789),.O(N789_NOT));
and2 gate( .a(N788_NOT), .b(p393), .O(EX981) );
and2 gate( .a(N789_NOT), .b(EX981), .O(EX982) );
and2 gate( .a(N788), .b(p394), .O(EX983) );
and2 gate( .a(N789_NOT), .b(EX983), .O(EX984) );
and2 gate( .a(N788_NOT), .b(p395), .O(EX985) );
and2 gate( .a(N789), .b(EX985), .O(EX986) );
and2 gate( .a(N788), .b(p396), .O(EX987) );
and2 gate( .a(N789), .b(EX987), .O(EX988) );
or2  gate( .a(EX982), .b(EX984), .O(EX989) );
or2  gate( .a(EX986), .b(EX989), .O(EX990) );
or2  gate( .a(EX988), .b(EX990), .O(N802) );
nor2 gate313( .a(N790), .b(N791), .O(N803) );
inv1 gate( .a(N792),.O(N792_NOT) );
inv1 gate( .a(N793),.O(N793_NOT));
and2 gate( .a(N792_NOT), .b(p397), .O(EX991) );
and2 gate( .a(N793_NOT), .b(EX991), .O(EX992) );
and2 gate( .a(N792), .b(p398), .O(EX993) );
and2 gate( .a(N793_NOT), .b(EX993), .O(EX994) );
and2 gate( .a(N792_NOT), .b(p399), .O(EX995) );
and2 gate( .a(N793), .b(EX995), .O(EX996) );
and2 gate( .a(N792), .b(p400), .O(EX997) );
and2 gate( .a(N793), .b(EX997), .O(EX998) );
or2  gate( .a(EX992), .b(EX994), .O(EX999) );
or2  gate( .a(EX996), .b(EX999), .O(EX1000) );
or2  gate( .a(EX998), .b(EX1000), .O(N804) );
inv1 gate( .a(N340),.O(N340_NOT) );
inv1 gate( .a(N794),.O(N794_NOT));
and2 gate( .a(N340_NOT), .b(p401), .O(EX1001) );
and2 gate( .a(N794_NOT), .b(EX1001), .O(EX1002) );
and2 gate( .a(N340), .b(p402), .O(EX1003) );
and2 gate( .a(N794_NOT), .b(EX1003), .O(EX1004) );
and2 gate( .a(N340_NOT), .b(p403), .O(EX1005) );
and2 gate( .a(N794), .b(EX1005), .O(EX1006) );
and2 gate( .a(N340), .b(p404), .O(EX1007) );
and2 gate( .a(N794), .b(EX1007), .O(EX1008) );
or2  gate( .a(EX1002), .b(EX1004), .O(EX1009) );
or2  gate( .a(EX1006), .b(EX1009), .O(EX1010) );
or2  gate( .a(EX1008), .b(EX1010), .O(N805) );
inv1 gate( .a(N692),.O(N692_NOT) );
inv1 gate( .a(N796),.O(N796_NOT));
and2 gate( .a(N692_NOT), .b(p405), .O(EX1011) );
and2 gate( .a(N796_NOT), .b(EX1011), .O(EX1012) );
and2 gate( .a(N692), .b(p406), .O(EX1013) );
and2 gate( .a(N796_NOT), .b(EX1013), .O(EX1014) );
and2 gate( .a(N692_NOT), .b(p407), .O(EX1015) );
and2 gate( .a(N796), .b(EX1015), .O(EX1016) );
and2 gate( .a(N692), .b(p408), .O(EX1017) );
and2 gate( .a(N796), .b(EX1017), .O(EX1018) );
or2  gate( .a(EX1012), .b(EX1014), .O(EX1019) );
or2  gate( .a(EX1016), .b(EX1019), .O(EX1020) );
or2  gate( .a(EX1018), .b(EX1020), .O(N806) );
inv1 gate( .a(N692),.O(N692_NOT) );
inv1 gate( .a(N796),.O(N796_NOT));
and2 gate( .a(N692_NOT), .b(p409), .O(EX1021) );
and2 gate( .a(N796_NOT), .b(EX1021), .O(EX1022) );
and2 gate( .a(N692), .b(p410), .O(EX1023) );
and2 gate( .a(N796_NOT), .b(EX1023), .O(EX1024) );
and2 gate( .a(N692_NOT), .b(p411), .O(EX1025) );
and2 gate( .a(N796), .b(EX1025), .O(EX1026) );
and2 gate( .a(N692), .b(p412), .O(EX1027) );
and2 gate( .a(N796), .b(EX1027), .O(EX1028) );
or2  gate( .a(EX1022), .b(EX1024), .O(EX1029) );
or2  gate( .a(EX1026), .b(EX1029), .O(EX1030) );
or2  gate( .a(EX1028), .b(EX1030), .O(N807) );
and2 gate318( .a(N219), .b(N802), .O(N808) );
and2 gate319( .a(N219), .b(N803), .O(N809) );
and2 gate320( .a(N219), .b(N804), .O(N810) );
nand4 gate321( .a(N805), .b(N787), .c(N731), .d(N529), .O(N811) );
nand2 gate322( .a(N619), .b(N796), .O(N812) );
nand3 gate323( .a(N609), .b(N619), .c(N796), .O(N813) );
nand4 gate324( .a(N600), .b(N609), .c(N619), .d(N796), .O(N814) );
nand4 gate325( .a(N738), .b(N765), .c(N766), .d(N814), .O(N815) );
nand3 gate326( .a(N741), .b(N764), .c(N813), .O(N819) );
nand2 gate327( .a(N744), .b(N812), .O(N822) );
nor2 gate328( .a(N806), .b(N807), .O(N825) );
inv1 gate( .a(N335),.O(N335_NOT) );
inv1 gate( .a(N808),.O(N808_NOT));
and2 gate( .a(N335_NOT), .b(p413), .O(EX1031) );
and2 gate( .a(N808_NOT), .b(EX1031), .O(EX1032) );
and2 gate( .a(N335), .b(p414), .O(EX1033) );
and2 gate( .a(N808_NOT), .b(EX1033), .O(EX1034) );
and2 gate( .a(N335_NOT), .b(p415), .O(EX1035) );
and2 gate( .a(N808), .b(EX1035), .O(EX1036) );
and2 gate( .a(N335), .b(p416), .O(EX1037) );
and2 gate( .a(N808), .b(EX1037), .O(EX1038) );
or2  gate( .a(EX1032), .b(EX1034), .O(EX1039) );
or2  gate( .a(EX1036), .b(EX1039), .O(EX1040) );
or2  gate( .a(EX1038), .b(EX1040), .O(N826) );
nor2 gate330( .a(N336), .b(N809), .O(N827) );
nor2 gate331( .a(N338), .b(N810), .O(N828) );
inv1 gate332( .a(N811), .O(N829) );
inv1 gate( .a(N665),.O(N665_NOT) );
inv1 gate( .a(N815),.O(N815_NOT));
and2 gate( .a(N665_NOT), .b(p417), .O(EX1041) );
and2 gate( .a(N815_NOT), .b(EX1041), .O(EX1042) );
and2 gate( .a(N665), .b(p418), .O(EX1043) );
and2 gate( .a(N815_NOT), .b(EX1043), .O(EX1044) );
and2 gate( .a(N665_NOT), .b(p419), .O(EX1045) );
and2 gate( .a(N815), .b(EX1045), .O(EX1046) );
and2 gate( .a(N665), .b(p420), .O(EX1047) );
and2 gate( .a(N815), .b(EX1047), .O(EX1048) );
or2  gate( .a(EX1042), .b(EX1044), .O(EX1049) );
or2  gate( .a(EX1046), .b(EX1049), .O(EX1050) );
or2  gate( .a(EX1048), .b(EX1050), .O(N830) );
inv1 gate( .a(N665),.O(N665_NOT) );
inv1 gate( .a(N815),.O(N815_NOT));
and2 gate( .a(N665_NOT), .b(p421), .O(EX1051) );
and2 gate( .a(N815_NOT), .b(EX1051), .O(EX1052) );
and2 gate( .a(N665), .b(p422), .O(EX1053) );
and2 gate( .a(N815_NOT), .b(EX1053), .O(EX1054) );
and2 gate( .a(N665_NOT), .b(p423), .O(EX1055) );
and2 gate( .a(N815), .b(EX1055), .O(EX1056) );
and2 gate( .a(N665), .b(p424), .O(EX1057) );
and2 gate( .a(N815), .b(EX1057), .O(EX1058) );
or2  gate( .a(EX1052), .b(EX1054), .O(EX1059) );
or2  gate( .a(EX1056), .b(EX1059), .O(EX1060) );
or2  gate( .a(EX1058), .b(EX1060), .O(N831) );
nor2 gate335( .a(N673), .b(N819), .O(N832) );
and2 gate336( .a(N673), .b(N819), .O(N833) );
nor2 gate337( .a(N682), .b(N822), .O(N834) );
inv1 gate( .a(N682),.O(N682_NOT) );
inv1 gate( .a(N822),.O(N822_NOT));
and2 gate( .a(N682_NOT), .b(p425), .O(EX1061) );
and2 gate( .a(N822_NOT), .b(EX1061), .O(EX1062) );
and2 gate( .a(N682), .b(p426), .O(EX1063) );
and2 gate( .a(N822_NOT), .b(EX1063), .O(EX1064) );
and2 gate( .a(N682_NOT), .b(p427), .O(EX1065) );
and2 gate( .a(N822), .b(EX1065), .O(EX1066) );
and2 gate( .a(N682), .b(p428), .O(EX1067) );
and2 gate( .a(N822), .b(EX1067), .O(EX1068) );
or2  gate( .a(EX1062), .b(EX1064), .O(EX1069) );
or2  gate( .a(EX1066), .b(EX1069), .O(EX1070) );
or2  gate( .a(EX1068), .b(EX1070), .O(N835) );
and2 gate339( .a(N219), .b(N825), .O(N836) );
nand3 gate340( .a(N826), .b(N777), .c(N704), .O(N837) );
nand4 gate341( .a(N827), .b(N781), .c(N712), .d(N527), .O(N838) );
nand4 gate342( .a(N828), .b(N785), .c(N721), .d(N528), .O(N839) );
inv1 gate343( .a(N829), .O(N840) );
inv1 gate( .a(N815),.O(N815_NOT) );
inv1 gate( .a(N593),.O(N593_NOT));
and2 gate( .a(N815_NOT), .b(p429), .O(EX1071) );
and2 gate( .a(N593_NOT), .b(EX1071), .O(EX1072) );
and2 gate( .a(N815), .b(p430), .O(EX1073) );
and2 gate( .a(N593_NOT), .b(EX1073), .O(EX1074) );
and2 gate( .a(N815_NOT), .b(p431), .O(EX1075) );
and2 gate( .a(N593), .b(EX1075), .O(EX1076) );
and2 gate( .a(N815), .b(p432), .O(EX1077) );
and2 gate( .a(N593), .b(EX1077), .O(EX1078) );
or2  gate( .a(EX1072), .b(EX1074), .O(EX1079) );
or2  gate( .a(EX1076), .b(EX1079), .O(EX1080) );
or2  gate( .a(EX1078), .b(EX1080), .O(N841) );
nor2 gate345( .a(N830), .b(N831), .O(N842) );
inv1 gate( .a(N832),.O(N832_NOT) );
inv1 gate( .a(N833),.O(N833_NOT));
and2 gate( .a(N832_NOT), .b(p433), .O(EX1081) );
and2 gate( .a(N833_NOT), .b(EX1081), .O(EX1082) );
and2 gate( .a(N832), .b(p434), .O(EX1083) );
and2 gate( .a(N833_NOT), .b(EX1083), .O(EX1084) );
and2 gate( .a(N832_NOT), .b(p435), .O(EX1085) );
and2 gate( .a(N833), .b(EX1085), .O(EX1086) );
and2 gate( .a(N832), .b(p436), .O(EX1087) );
and2 gate( .a(N833), .b(EX1087), .O(EX1088) );
or2  gate( .a(EX1082), .b(EX1084), .O(EX1089) );
or2  gate( .a(EX1086), .b(EX1089), .O(EX1090) );
or2  gate( .a(EX1088), .b(EX1090), .O(N843) );
nor2 gate347( .a(N834), .b(N835), .O(N844) );
nor2 gate348( .a(N334), .b(N836), .O(N845) );
inv1 gate349( .a(N837), .O(N846) );
inv1 gate350( .a(N838), .O(N847) );
inv1 gate351( .a(N839), .O(N848) );
and2 gate352( .a(N735), .b(N841), .O(N849) );
buf1 gate353( .a(N840), .O(N850) );
inv1 gate( .a(N219),.O(N219_NOT) );
inv1 gate( .a(N842),.O(N842_NOT));
and2 gate( .a(N219_NOT), .b(p437), .O(EX1091) );
and2 gate( .a(N842_NOT), .b(EX1091), .O(EX1092) );
and2 gate( .a(N219), .b(p438), .O(EX1093) );
and2 gate( .a(N842_NOT), .b(EX1093), .O(EX1094) );
and2 gate( .a(N219_NOT), .b(p439), .O(EX1095) );
and2 gate( .a(N842), .b(EX1095), .O(EX1096) );
and2 gate( .a(N219), .b(p440), .O(EX1097) );
and2 gate( .a(N842), .b(EX1097), .O(EX1098) );
or2  gate( .a(EX1092), .b(EX1094), .O(EX1099) );
or2  gate( .a(EX1096), .b(EX1099), .O(EX1100) );
or2  gate( .a(EX1098), .b(EX1100), .O(N851) );
and2 gate355( .a(N219), .b(N843), .O(N852) );
and2 gate356( .a(N219), .b(N844), .O(N853) );
nand3 gate357( .a(N845), .b(N772), .c(N696), .O(N854) );
inv1 gate358( .a(N846), .O(N855) );
inv1 gate359( .a(N847), .O(N856) );
inv1 gate360( .a(N848), .O(N857) );
inv1 gate361( .a(N849), .O(N858) );
inv1 gate( .a(N417),.O(N417_NOT) );
inv1 gate( .a(N851),.O(N851_NOT));
and2 gate( .a(N417_NOT), .b(p441), .O(EX1101) );
and2 gate( .a(N851_NOT), .b(EX1101), .O(EX1102) );
and2 gate( .a(N417), .b(p442), .O(EX1103) );
and2 gate( .a(N851_NOT), .b(EX1103), .O(EX1104) );
and2 gate( .a(N417_NOT), .b(p443), .O(EX1105) );
and2 gate( .a(N851), .b(EX1105), .O(EX1106) );
and2 gate( .a(N417), .b(p444), .O(EX1107) );
and2 gate( .a(N851), .b(EX1107), .O(EX1108) );
or2  gate( .a(EX1102), .b(EX1104), .O(EX1109) );
or2  gate( .a(EX1106), .b(EX1109), .O(EX1110) );
or2  gate( .a(EX1108), .b(EX1110), .O(N859) );
nor2 gate363( .a(N332), .b(N852), .O(N860) );
nor2 gate364( .a(N333), .b(N853), .O(N861) );
inv1 gate365( .a(N854), .O(N862) );
buf1 gate366( .a(N855), .O(N863) );
buf1 gate367( .a(N856), .O(N864) );
buf1 gate368( .a(N857), .O(N865) );
buf1 gate369( .a(N858), .O(N866) );
nand3 gate370( .a(N859), .b(N769), .c(N669), .O(N867) );
nand3 gate371( .a(N860), .b(N770), .c(N677), .O(N868) );
nand3 gate372( .a(N861), .b(N771), .c(N686), .O(N869) );
inv1 gate373( .a(N862), .O(N870) );
inv1 gate374( .a(N867), .O(N871) );
inv1 gate375( .a(N868), .O(N872) );
inv1 gate376( .a(N869), .O(N873) );
buf1 gate377( .a(N870), .O(N874) );
inv1 gate378( .a(N871), .O(N875) );
inv1 gate379( .a(N872), .O(N876) );
inv1 gate380( .a(N873), .O(N877) );
buf1 gate381( .a(N875), .O(N878) );
buf1 gate382( .a(N876), .O(N879) );
buf1 gate383( .a(N877), .O(N880) );

endmodule
