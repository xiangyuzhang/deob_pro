
module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;

input p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,
        p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,
        p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,
        p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,
        p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,
        p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,
        p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,
        p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,
        p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,
        p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,
        p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,
        p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,
        p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,
        p131,p132;

output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429,
     N118_NOT,N4_NOT,N8_NOT,N119_NOT,N130_NOT,N43_NOT,N138_NOT,N69_NOT,N142_NOT,N82_NOT,
     N150_NOT,N108_NOT,N27_NOT,N123_NOT,N66_NOT,N135_NOT,N73_NOT,N139_NOT,N79_NOT,N139_NOT,
     N112_NOT,N151_NOT,N115_NOT,N151_NOT,N203_NOT,N165_NOT,N203_NOT,N171_NOT,N203_NOT,N174_NOT,
     N203_NOT,N180_NOT,N213_NOT,N37_NOT,N213_NOT,N89_NOT,N213_NOT,N102_NOT,N239_NOT,N191_NOT,
     N243_NOT,N193_NOT,N251_NOT,N197_NOT,N230_NOT,N186_NOT,N233_NOT,N188_NOT,N236_NOT,N190_NOT,
     N247_NOT,N196_NOT,N309_NOT,N267_NOT,N309_NOT,N276_NOT,N319_NOT,N34_NOT,N343_NOT,N308_NOT,
     N360_NOT,N27_NOT,N360_NOT,N66_NOT,N360_NOT,N105_NOT,EX1,EX2,EX3,EX4,EX5,EX6,EX7,EX8,EX9,EX10,
     EX11,EX12,EX13,EX14,EX15,EX16,EX17,EX18,EX19,EX20,
     EX21,EX22,EX23,EX24,EX25,EX26,EX27,EX28,EX29,EX30,
     EX31,EX32,EX33,EX34,EX35,EX36,EX37,EX38,EX39,EX40,
     EX41,EX42,EX43,EX44,EX45,EX46,EX47,EX48,EX49,EX50,
     EX51,EX52,EX53,EX54,EX55,EX56,EX57,EX58,EX59,EX60,
     EX61,EX62,EX63,EX64,EX65,EX66,EX67,EX68,EX69,EX70,
     EX71,EX72,EX73,EX74,EX75,EX76,EX77,EX78,EX79,EX80,
     EX81,EX82,EX83,EX84,EX85,EX86,EX87,EX88,EX89,EX90,
     EX91,EX92,EX93,EX94,EX95,EX96,EX97,EX98,EX99,EX100,
     EX101,EX102,EX103,EX104,EX105,EX106,EX107,EX108,EX109,EX110,
     EX111,EX112,EX113,EX114,EX115,EX116,EX117,EX118,EX119,EX120,
     EX121,EX122,EX123,EX124,EX125,EX126,EX127,EX128,EX129,EX130,
     EX131,EX132,EX133,EX134,EX135,EX136,EX137,EX138,EX139,EX140,
     EX141,EX142,EX143,EX144,EX145,EX146,EX147,EX148,EX149,EX150,
     EX151,EX152,EX153,EX154,EX155,EX156,EX157,EX158,EX159,EX160,
     EX161,EX162,EX163,EX164,EX165,EX166,EX167,EX168,EX169,EX170,
     EX171,EX172,EX173,EX174,EX175,EX176,EX177,EX178,EX179,EX180,
     EX181,EX182,EX183,EX184,EX185,EX186,EX187,EX188,EX189,EX190,
     EX191,EX192,EX193,EX194,EX195,EX196,EX197,EX198,EX199,EX200,
     EX201,EX202,EX203,EX204,EX205,EX206,EX207,EX208,EX209,EX210,
     EX211,EX212,EX213,EX214,EX215,EX216,EX217,EX218,EX219,EX220,
     EX221,EX222,EX223,EX224,EX225,EX226,EX227,EX228,EX229,EX230,
     EX231,EX232,EX233,EX234,EX235,EX236,EX237,EX238,EX239,EX240,
     EX241,EX242,EX243,EX244,EX245,EX246,EX247,EX248,EX249,EX250,
     EX251,EX252,EX253,EX254,EX255,EX256,EX257,EX258,EX259,EX260,
     EX261,EX262,EX263,EX264,EX265,EX266,EX267,EX268,EX269,EX270,
     EX271,EX272,EX273,EX274,EX275,EX276,EX277,EX278,EX279,EX280,
     EX281,EX282,EX283,EX284,EX285,EX286,EX287,EX288,EX289,EX290,
     EX291,EX292,EX293,EX294,EX295,EX296,EX297,EX298,EX299,EX300,
     EX301,EX302,EX303,EX304,EX305,EX306,EX307,EX308,EX309,EX310,
     EX311,EX312,EX313,EX314,EX315,EX316,EX317,EX318,EX319,EX320,
     EX321,EX322,EX323,EX324,EX325,EX326,EX327,EX328,EX329,EX330;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
inv1 gate( .a(N118),.O(N118_NOT) );
inv1 gate( .a(N4),.O(N4_NOT));
and2 gate( .a(N118_NOT), .b(p1), .O(EX1) );
and2 gate( .a(N4_NOT), .b(EX1), .O(EX2) );
and2 gate( .a(N118), .b(p2), .O(EX3) );
and2 gate( .a(N4_NOT), .b(EX3), .O(EX4) );
and2 gate( .a(N118_NOT), .b(p3), .O(EX5) );
and2 gate( .a(N4), .b(EX5), .O(EX6) );
and2 gate( .a(N118), .b(p4), .O(EX7) );
and2 gate( .a(N4), .b(EX7), .O(EX8) );
or2  gate( .a(EX2), .b(EX4), .O(EX9) );
or2  gate( .a(EX6), .b(EX9), .O(EX10) );
or2  gate( .a(EX8), .b(EX10), .O(N154) );
inv1 gate( .a(N8),.O(N8_NOT) );
inv1 gate( .a(N119),.O(N119_NOT));
and2 gate( .a(N8_NOT), .b(p5), .O(EX11) );
and2 gate( .a(N119_NOT), .b(EX11), .O(EX12) );
and2 gate( .a(N8), .b(p6), .O(EX13) );
and2 gate( .a(N119_NOT), .b(EX13), .O(EX14) );
and2 gate( .a(N8_NOT), .b(p7), .O(EX15) );
and2 gate( .a(N119), .b(EX15), .O(EX16) );
and2 gate( .a(N8), .b(p8), .O(EX17) );
and2 gate( .a(N119), .b(EX17), .O(EX18) );
or2  gate( .a(EX12), .b(EX14), .O(EX19) );
or2  gate( .a(EX16), .b(EX19), .O(EX20) );
or2  gate( .a(EX18), .b(EX20), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );
nand2 gate23( .a(N126), .b(N30), .O(N162) );
inv1 gate( .a(N130),.O(N130_NOT) );
inv1 gate( .a(N43),.O(N43_NOT));
and2 gate( .a(N130_NOT), .b(p9), .O(EX21) );
and2 gate( .a(N43_NOT), .b(EX21), .O(EX22) );
and2 gate( .a(N130), .b(p10), .O(EX23) );
and2 gate( .a(N43_NOT), .b(EX23), .O(EX24) );
and2 gate( .a(N130_NOT), .b(p11), .O(EX25) );
and2 gate( .a(N43), .b(EX25), .O(EX26) );
and2 gate( .a(N130), .b(p12), .O(EX27) );
and2 gate( .a(N43), .b(EX27), .O(EX28) );
or2  gate( .a(EX22), .b(EX24), .O(EX29) );
or2  gate( .a(EX26), .b(EX29), .O(EX30) );
or2  gate( .a(EX28), .b(EX30), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );
inv1 gate( .a(N138),.O(N138_NOT) );
inv1 gate( .a(N69),.O(N69_NOT));
and2 gate( .a(N138_NOT), .b(p13), .O(EX31) );
and2 gate( .a(N69_NOT), .b(EX31), .O(EX32) );
and2 gate( .a(N138), .b(p14), .O(EX33) );
and2 gate( .a(N69_NOT), .b(EX33), .O(EX34) );
and2 gate( .a(N138_NOT), .b(p15), .O(EX35) );
and2 gate( .a(N69), .b(EX35), .O(EX36) );
and2 gate( .a(N138), .b(p16), .O(EX37) );
and2 gate( .a(N69), .b(EX37), .O(EX38) );
or2  gate( .a(EX32), .b(EX34), .O(EX39) );
or2  gate( .a(EX36), .b(EX39), .O(EX40) );
or2  gate( .a(EX38), .b(EX40), .O(N171) );
inv1 gate( .a(N142),.O(N142_NOT) );
inv1 gate( .a(N82),.O(N82_NOT));
and2 gate( .a(N142_NOT), .b(p17), .O(EX41) );
and2 gate( .a(N82_NOT), .b(EX41), .O(EX42) );
and2 gate( .a(N142), .b(p18), .O(EX43) );
and2 gate( .a(N82_NOT), .b(EX43), .O(EX44) );
and2 gate( .a(N142_NOT), .b(p19), .O(EX45) );
and2 gate( .a(N82), .b(EX45), .O(EX46) );
and2 gate( .a(N142), .b(p20), .O(EX47) );
and2 gate( .a(N82), .b(EX47), .O(EX48) );
or2  gate( .a(EX42), .b(EX44), .O(EX49) );
or2  gate( .a(EX46), .b(EX49), .O(EX50) );
or2  gate( .a(EX48), .b(EX50), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );
inv1 gate( .a(N150),.O(N150_NOT) );
inv1 gate( .a(N108),.O(N108_NOT));
and2 gate( .a(N150_NOT), .b(p21), .O(EX51) );
and2 gate( .a(N108_NOT), .b(EX51), .O(EX52) );
and2 gate( .a(N150), .b(p22), .O(EX53) );
and2 gate( .a(N108_NOT), .b(EX53), .O(EX54) );
and2 gate( .a(N150_NOT), .b(p23), .O(EX55) );
and2 gate( .a(N108), .b(EX55), .O(EX56) );
and2 gate( .a(N150), .b(p24), .O(EX57) );
and2 gate( .a(N108), .b(EX57), .O(EX58) );
or2  gate( .a(EX52), .b(EX54), .O(EX59) );
or2  gate( .a(EX56), .b(EX59), .O(EX60) );
or2  gate( .a(EX58), .b(EX60), .O(N180) );
nor2 gate30( .a(N21), .b(N123), .O(N183) );
inv1 gate( .a(N27),.O(N27_NOT) );
inv1 gate( .a(N123),.O(N123_NOT));
and2 gate( .a(N27_NOT), .b(p25), .O(EX61) );
and2 gate( .a(N123_NOT), .b(EX61), .O(EX62) );
and2 gate( .a(N27), .b(p26), .O(EX63) );
and2 gate( .a(N123_NOT), .b(EX63), .O(EX64) );
and2 gate( .a(N27_NOT), .b(p27), .O(EX65) );
and2 gate( .a(N123), .b(EX65), .O(EX66) );
and2 gate( .a(N27), .b(p28), .O(EX67) );
and2 gate( .a(N123), .b(EX67), .O(EX68) );
or2  gate( .a(EX62), .b(EX64), .O(EX69) );
or2  gate( .a(EX66), .b(EX69), .O(EX70) );
or2  gate( .a(EX68), .b(EX70), .O(N184) );
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );
nor2 gate36( .a(N60), .b(N135), .O(N189) );
inv1 gate( .a(N66),.O(N66_NOT) );
inv1 gate( .a(N135),.O(N135_NOT));
and2 gate( .a(N66_NOT), .b(p29), .O(EX71) );
and2 gate( .a(N135_NOT), .b(EX71), .O(EX72) );
and2 gate( .a(N66), .b(p30), .O(EX73) );
and2 gate( .a(N135_NOT), .b(EX73), .O(EX74) );
and2 gate( .a(N66_NOT), .b(p31), .O(EX75) );
and2 gate( .a(N135), .b(EX75), .O(EX76) );
and2 gate( .a(N66), .b(p32), .O(EX77) );
and2 gate( .a(N135), .b(EX77), .O(EX78) );
or2  gate( .a(EX72), .b(EX74), .O(EX79) );
or2  gate( .a(EX76), .b(EX79), .O(EX80) );
or2  gate( .a(EX78), .b(EX80), .O(N190) );
inv1 gate( .a(N73),.O(N73_NOT) );
inv1 gate( .a(N139),.O(N139_NOT));
and2 gate( .a(N73_NOT), .b(p33), .O(EX81) );
and2 gate( .a(N139_NOT), .b(EX81), .O(EX82) );
and2 gate( .a(N73), .b(p34), .O(EX83) );
and2 gate( .a(N139_NOT), .b(EX83), .O(EX84) );
and2 gate( .a(N73_NOT), .b(p35), .O(EX85) );
and2 gate( .a(N139), .b(EX85), .O(EX86) );
and2 gate( .a(N73), .b(p36), .O(EX87) );
and2 gate( .a(N139), .b(EX87), .O(EX88) );
or2  gate( .a(EX82), .b(EX84), .O(EX89) );
or2  gate( .a(EX86), .b(EX89), .O(EX90) );
or2  gate( .a(EX88), .b(EX90), .O(N191) );
inv1 gate( .a(N79),.O(N79_NOT) );
inv1 gate( .a(N139),.O(N139_NOT));
and2 gate( .a(N79_NOT), .b(p37), .O(EX91) );
and2 gate( .a(N139_NOT), .b(EX91), .O(EX92) );
and2 gate( .a(N79), .b(p38), .O(EX93) );
and2 gate( .a(N139_NOT), .b(EX93), .O(EX94) );
and2 gate( .a(N79_NOT), .b(p39), .O(EX95) );
and2 gate( .a(N139), .b(EX95), .O(EX96) );
and2 gate( .a(N79), .b(p40), .O(EX97) );
and2 gate( .a(N139), .b(EX97), .O(EX98) );
or2  gate( .a(EX92), .b(EX94), .O(EX99) );
or2  gate( .a(EX96), .b(EX99), .O(EX100) );
or2  gate( .a(EX98), .b(EX100), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );
nor2 gate41( .a(N92), .b(N143), .O(N194) );
nor2 gate42( .a(N99), .b(N147), .O(N195) );
nor2 gate43( .a(N105), .b(N147), .O(N196) );
inv1 gate( .a(N112),.O(N112_NOT) );
inv1 gate( .a(N151),.O(N151_NOT));
and2 gate( .a(N112_NOT), .b(p41), .O(EX101) );
and2 gate( .a(N151_NOT), .b(EX101), .O(EX102) );
and2 gate( .a(N112), .b(p42), .O(EX103) );
and2 gate( .a(N151_NOT), .b(EX103), .O(EX104) );
and2 gate( .a(N112_NOT), .b(p43), .O(EX105) );
and2 gate( .a(N151), .b(EX105), .O(EX106) );
and2 gate( .a(N112), .b(p44), .O(EX107) );
and2 gate( .a(N151), .b(EX107), .O(EX108) );
or2  gate( .a(EX102), .b(EX104), .O(EX109) );
or2  gate( .a(EX106), .b(EX109), .O(EX110) );
or2  gate( .a(EX108), .b(EX110), .O(N197) );
inv1 gate( .a(N115),.O(N115_NOT) );
inv1 gate( .a(N151),.O(N151_NOT));
and2 gate( .a(N115_NOT), .b(p45), .O(EX111) );
and2 gate( .a(N151_NOT), .b(EX111), .O(EX112) );
and2 gate( .a(N115), .b(p46), .O(EX113) );
and2 gate( .a(N151_NOT), .b(EX113), .O(EX114) );
and2 gate( .a(N115_NOT), .b(p47), .O(EX115) );
and2 gate( .a(N151), .b(EX115), .O(EX116) );
and2 gate( .a(N115), .b(p48), .O(EX117) );
and2 gate( .a(N151), .b(EX117), .O(EX118) );
or2  gate( .a(EX112), .b(EX114), .O(EX119) );
or2  gate( .a(EX116), .b(EX119), .O(EX120) );
or2  gate( .a(EX118), .b(EX120), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );
xor2 gate52( .a(N203), .b(N162), .O(N230) );
inv1 gate( .a(N203),.O(N203_NOT) );
inv1 gate( .a(N165),.O(N165_NOT));
and2 gate( .a(N203_NOT), .b(p49), .O(EX121) );
and2 gate( .a(N165_NOT), .b(EX121), .O(EX122) );
and2 gate( .a(N203), .b(p50), .O(EX123) );
and2 gate( .a(N165_NOT), .b(EX123), .O(EX124) );
and2 gate( .a(N203_NOT), .b(p51), .O(EX125) );
and2 gate( .a(N165), .b(EX125), .O(EX126) );
and2 gate( .a(N203), .b(p52), .O(EX127) );
and2 gate( .a(N165), .b(EX127), .O(EX128) );
or2  gate( .a(EX122), .b(EX124), .O(EX129) );
or2  gate( .a(EX126), .b(EX129), .O(EX130) );
or2  gate( .a(EX128), .b(EX130), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );
inv1 gate( .a(N203),.O(N203_NOT) );
inv1 gate( .a(N171),.O(N171_NOT));
and2 gate( .a(N203_NOT), .b(p53), .O(EX131) );
and2 gate( .a(N171_NOT), .b(EX131), .O(EX132) );
and2 gate( .a(N203), .b(p54), .O(EX133) );
and2 gate( .a(N171_NOT), .b(EX133), .O(EX134) );
and2 gate( .a(N203_NOT), .b(p55), .O(EX135) );
and2 gate( .a(N171), .b(EX135), .O(EX136) );
and2 gate( .a(N203), .b(p56), .O(EX137) );
and2 gate( .a(N171), .b(EX137), .O(EX138) );
or2  gate( .a(EX132), .b(EX134), .O(EX139) );
or2  gate( .a(EX136), .b(EX139), .O(EX140) );
or2  gate( .a(EX138), .b(EX140), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );
inv1 gate( .a(N203),.O(N203_NOT) );
inv1 gate( .a(N174),.O(N174_NOT));
and2 gate( .a(N203_NOT), .b(p57), .O(EX141) );
and2 gate( .a(N174_NOT), .b(EX141), .O(EX142) );
and2 gate( .a(N203), .b(p58), .O(EX143) );
and2 gate( .a(N174_NOT), .b(EX143), .O(EX144) );
and2 gate( .a(N203_NOT), .b(p59), .O(EX145) );
and2 gate( .a(N174), .b(EX145), .O(EX146) );
and2 gate( .a(N203), .b(p60), .O(EX147) );
and2 gate( .a(N174), .b(EX147), .O(EX148) );
or2  gate( .a(EX142), .b(EX144), .O(EX149) );
or2  gate( .a(EX146), .b(EX149), .O(EX150) );
or2  gate( .a(EX148), .b(EX150), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24), .O(N250) );
inv1 gate( .a(N203),.O(N203_NOT) );
inv1 gate( .a(N180),.O(N180_NOT));
and2 gate( .a(N203_NOT), .b(p61), .O(EX151) );
and2 gate( .a(N180_NOT), .b(EX151), .O(EX152) );
and2 gate( .a(N203), .b(p62), .O(EX153) );
and2 gate( .a(N180_NOT), .b(EX153), .O(EX154) );
and2 gate( .a(N203_NOT), .b(p63), .O(EX155) );
and2 gate( .a(N180), .b(EX155), .O(EX156) );
and2 gate( .a(N203), .b(p64), .O(EX157) );
and2 gate( .a(N180), .b(EX157), .O(EX158) );
or2  gate( .a(EX152), .b(EX154), .O(EX159) );
or2  gate( .a(EX156), .b(EX159), .O(EX160) );
or2  gate( .a(EX158), .b(EX160), .O(N251) );
inv1 gate( .a(N213),.O(N213_NOT) );
inv1 gate( .a(N37),.O(N37_NOT));
and2 gate( .a(N213_NOT), .b(p65), .O(EX161) );
and2 gate( .a(N37_NOT), .b(EX161), .O(EX162) );
and2 gate( .a(N213), .b(p66), .O(EX163) );
and2 gate( .a(N37_NOT), .b(EX163), .O(EX164) );
and2 gate( .a(N213_NOT), .b(p67), .O(EX165) );
and2 gate( .a(N37), .b(EX165), .O(EX166) );
and2 gate( .a(N213), .b(p68), .O(EX167) );
and2 gate( .a(N37), .b(EX167), .O(EX168) );
or2  gate( .a(EX162), .b(EX164), .O(EX169) );
or2  gate( .a(EX166), .b(EX169), .O(EX170) );
or2  gate( .a(EX168), .b(EX170), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );
inv1 gate( .a(N213),.O(N213_NOT) );
inv1 gate( .a(N89),.O(N89_NOT));
and2 gate( .a(N213_NOT), .b(p69), .O(EX171) );
and2 gate( .a(N89_NOT), .b(EX171), .O(EX172) );
and2 gate( .a(N213), .b(p70), .O(EX173) );
and2 gate( .a(N89_NOT), .b(EX173), .O(EX174) );
and2 gate( .a(N213_NOT), .b(p71), .O(EX175) );
and2 gate( .a(N89), .b(EX175), .O(EX176) );
and2 gate( .a(N213), .b(p72), .O(EX177) );
and2 gate( .a(N89), .b(EX177), .O(EX178) );
or2  gate( .a(EX172), .b(EX174), .O(EX179) );
or2  gate( .a(EX176), .b(EX179), .O(EX180) );
or2  gate( .a(EX178), .b(EX180), .O(N258) );
inv1 gate( .a(N213),.O(N213_NOT) );
inv1 gate( .a(N102),.O(N102_NOT));
and2 gate( .a(N213_NOT), .b(p73), .O(EX181) );
and2 gate( .a(N102_NOT), .b(EX181), .O(EX182) );
and2 gate( .a(N213), .b(p74), .O(EX183) );
and2 gate( .a(N102_NOT), .b(EX183), .O(EX184) );
and2 gate( .a(N213_NOT), .b(p75), .O(EX185) );
and2 gate( .a(N102), .b(EX185), .O(EX186) );
and2 gate( .a(N213), .b(p76), .O(EX187) );
and2 gate( .a(N102), .b(EX187), .O(EX188) );
or2  gate( .a(EX182), .b(EX184), .O(EX189) );
or2  gate( .a(EX186), .b(EX189), .O(EX190) );
or2  gate( .a(EX188), .b(EX190), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );
nand2 gate71( .a(N230), .b(N185), .O(N267) );
nand2 gate72( .a(N233), .b(N187), .O(N270) );
nand2 gate73( .a(N236), .b(N189), .O(N273) );
inv1 gate( .a(N239),.O(N239_NOT) );
inv1 gate( .a(N191),.O(N191_NOT));
and2 gate( .a(N239_NOT), .b(p77), .O(EX191) );
and2 gate( .a(N191_NOT), .b(EX191), .O(EX192) );
and2 gate( .a(N239), .b(p78), .O(EX193) );
and2 gate( .a(N191_NOT), .b(EX193), .O(EX194) );
and2 gate( .a(N239_NOT), .b(p79), .O(EX195) );
and2 gate( .a(N191), .b(EX195), .O(EX196) );
and2 gate( .a(N239), .b(p80), .O(EX197) );
and2 gate( .a(N191), .b(EX197), .O(EX198) );
or2  gate( .a(EX192), .b(EX194), .O(EX199) );
or2  gate( .a(EX196), .b(EX199), .O(EX200) );
or2  gate( .a(EX198), .b(EX200), .O(N276) );
inv1 gate( .a(N243),.O(N243_NOT) );
inv1 gate( .a(N193),.O(N193_NOT));
and2 gate( .a(N243_NOT), .b(p81), .O(EX201) );
and2 gate( .a(N193_NOT), .b(EX201), .O(EX202) );
and2 gate( .a(N243), .b(p82), .O(EX203) );
and2 gate( .a(N193_NOT), .b(EX203), .O(EX204) );
and2 gate( .a(N243_NOT), .b(p83), .O(EX205) );
and2 gate( .a(N193), .b(EX205), .O(EX206) );
and2 gate( .a(N243), .b(p84), .O(EX207) );
and2 gate( .a(N193), .b(EX207), .O(EX208) );
or2  gate( .a(EX202), .b(EX204), .O(EX209) );
or2  gate( .a(EX206), .b(EX209), .O(EX210) );
or2  gate( .a(EX208), .b(EX210), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );
inv1 gate( .a(N251),.O(N251_NOT) );
inv1 gate( .a(N197),.O(N197_NOT));
and2 gate( .a(N251_NOT), .b(p85), .O(EX211) );
and2 gate( .a(N197_NOT), .b(EX211), .O(EX212) );
and2 gate( .a(N251), .b(p86), .O(EX213) );
and2 gate( .a(N197_NOT), .b(EX213), .O(EX214) );
and2 gate( .a(N251_NOT), .b(p87), .O(EX215) );
and2 gate( .a(N197), .b(EX215), .O(EX216) );
and2 gate( .a(N251), .b(p88), .O(EX217) );
and2 gate( .a(N197), .b(EX217), .O(EX218) );
or2  gate( .a(EX212), .b(EX214), .O(EX219) );
or2  gate( .a(EX216), .b(EX219), .O(EX220) );
or2  gate( .a(EX218), .b(EX220), .O(N285) );
nand2 gate78( .a(N227), .b(N184), .O(N288) );
inv1 gate( .a(N230),.O(N230_NOT) );
inv1 gate( .a(N186),.O(N186_NOT));
and2 gate( .a(N230_NOT), .b(p89), .O(EX221) );
and2 gate( .a(N186_NOT), .b(EX221), .O(EX222) );
and2 gate( .a(N230), .b(p90), .O(EX223) );
and2 gate( .a(N186_NOT), .b(EX223), .O(EX224) );
and2 gate( .a(N230_NOT), .b(p91), .O(EX225) );
and2 gate( .a(N186), .b(EX225), .O(EX226) );
and2 gate( .a(N230), .b(p92), .O(EX227) );
and2 gate( .a(N186), .b(EX227), .O(EX228) );
or2  gate( .a(EX222), .b(EX224), .O(EX229) );
or2  gate( .a(EX226), .b(EX229), .O(EX230) );
or2  gate( .a(EX228), .b(EX230), .O(N289) );
inv1 gate( .a(N233),.O(N233_NOT) );
inv1 gate( .a(N188),.O(N188_NOT));
and2 gate( .a(N233_NOT), .b(p93), .O(EX231) );
and2 gate( .a(N188_NOT), .b(EX231), .O(EX232) );
and2 gate( .a(N233), .b(p94), .O(EX233) );
and2 gate( .a(N188_NOT), .b(EX233), .O(EX234) );
and2 gate( .a(N233_NOT), .b(p95), .O(EX235) );
and2 gate( .a(N188), .b(EX235), .O(EX236) );
and2 gate( .a(N233), .b(p96), .O(EX237) );
and2 gate( .a(N188), .b(EX237), .O(EX238) );
or2  gate( .a(EX232), .b(EX234), .O(EX239) );
or2  gate( .a(EX236), .b(EX239), .O(EX240) );
or2  gate( .a(EX238), .b(EX240), .O(N290) );
inv1 gate( .a(N236),.O(N236_NOT) );
inv1 gate( .a(N190),.O(N190_NOT));
and2 gate( .a(N236_NOT), .b(p97), .O(EX241) );
and2 gate( .a(N190_NOT), .b(EX241), .O(EX242) );
and2 gate( .a(N236), .b(p98), .O(EX243) );
and2 gate( .a(N190_NOT), .b(EX243), .O(EX244) );
and2 gate( .a(N236_NOT), .b(p99), .O(EX245) );
and2 gate( .a(N190), .b(EX245), .O(EX246) );
and2 gate( .a(N236), .b(p100), .O(EX247) );
and2 gate( .a(N190), .b(EX247), .O(EX248) );
or2  gate( .a(EX242), .b(EX244), .O(EX249) );
or2  gate( .a(EX246), .b(EX249), .O(EX250) );
or2  gate( .a(EX248), .b(EX250), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );
inv1 gate( .a(N247),.O(N247_NOT) );
inv1 gate( .a(N196),.O(N196_NOT));
and2 gate( .a(N247_NOT), .b(p101), .O(EX251) );
and2 gate( .a(N196_NOT), .b(EX251), .O(EX252) );
and2 gate( .a(N247), .b(p102), .O(EX253) );
and2 gate( .a(N196_NOT), .b(EX253), .O(EX254) );
and2 gate( .a(N247_NOT), .b(p103), .O(EX255) );
and2 gate( .a(N196), .b(EX255), .O(EX256) );
and2 gate( .a(N247), .b(p104), .O(EX257) );
and2 gate( .a(N196), .b(EX257), .O(EX258) );
or2  gate( .a(EX252), .b(EX254), .O(EX259) );
or2  gate( .a(EX256), .b(EX259), .O(EX260) );
or2  gate( .a(EX258), .b(EX260), .O(N294) );
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );
inv1 gate( .a(N309),.O(N309_NOT) );
inv1 gate( .a(N267),.O(N267_NOT));
and2 gate( .a(N309_NOT), .b(p105), .O(EX261) );
and2 gate( .a(N267_NOT), .b(EX261), .O(EX262) );
and2 gate( .a(N309), .b(p106), .O(EX263) );
and2 gate( .a(N267_NOT), .b(EX263), .O(EX264) );
and2 gate( .a(N309_NOT), .b(p107), .O(EX265) );
and2 gate( .a(N267), .b(EX265), .O(EX266) );
and2 gate( .a(N309), .b(p108), .O(EX267) );
and2 gate( .a(N267), .b(EX267), .O(EX268) );
or2  gate( .a(EX262), .b(EX264), .O(EX269) );
or2  gate( .a(EX266), .b(EX269), .O(EX270) );
or2  gate( .a(EX268), .b(EX270), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );
inv1 gate( .a(N309),.O(N309_NOT) );
inv1 gate( .a(N276),.O(N276_NOT));
and2 gate( .a(N309_NOT), .b(p109), .O(EX271) );
and2 gate( .a(N276_NOT), .b(EX271), .O(EX272) );
and2 gate( .a(N309), .b(p110), .O(EX273) );
and2 gate( .a(N276_NOT), .b(EX273), .O(EX274) );
and2 gate( .a(N309_NOT), .b(p111), .O(EX275) );
and2 gate( .a(N276), .b(EX275), .O(EX276) );
and2 gate( .a(N309), .b(p112), .O(EX277) );
and2 gate( .a(N276), .b(EX277), .O(EX278) );
or2  gate( .a(EX272), .b(EX274), .O(EX279) );
or2  gate( .a(EX276), .b(EX279), .O(EX280) );
or2  gate( .a(EX278), .b(EX280), .O(N337) );
inv1 gate( .a(N319),.O(N319_NOT) );
inv1 gate( .a(N34),.O(N34_NOT));
and2 gate( .a(N319_NOT), .b(p113), .O(EX281) );
and2 gate( .a(N34_NOT), .b(EX281), .O(EX282) );
and2 gate( .a(N319), .b(p114), .O(EX283) );
and2 gate( .a(N34_NOT), .b(EX283), .O(EX284) );
and2 gate( .a(N319_NOT), .b(p115), .O(EX285) );
and2 gate( .a(N34), .b(EX285), .O(EX286) );
and2 gate( .a(N319), .b(p116), .O(EX287) );
and2 gate( .a(N34), .b(EX287), .O(EX288) );
or2  gate( .a(EX282), .b(EX284), .O(EX289) );
or2  gate( .a(EX286), .b(EX289), .O(EX290) );
or2  gate( .a(EX288), .b(EX290), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );
nand2 gate111( .a(N319), .b(N60), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );
nand2 gate113( .a(N319), .b(N73), .O(N344) );
nand2 gate114( .a(N319), .b(N86), .O(N345) );
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302), .O(N350) );
nand2 gate120( .a(N333), .b(N303), .O(N351) );
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );
inv1 gate( .a(N343),.O(N343_NOT) );
inv1 gate( .a(N308),.O(N308_NOT));
and2 gate( .a(N343_NOT), .b(p117), .O(EX291) );
and2 gate( .a(N308_NOT), .b(EX291), .O(EX292) );
and2 gate( .a(N343), .b(p118), .O(EX293) );
and2 gate( .a(N308_NOT), .b(EX293), .O(EX294) );
and2 gate( .a(N343_NOT), .b(p119), .O(EX295) );
and2 gate( .a(N308), .b(EX295), .O(EX296) );
and2 gate( .a(N343), .b(p120), .O(EX297) );
and2 gate( .a(N308), .b(EX297), .O(EX298) );
or2  gate( .a(EX292), .b(EX294), .O(EX299) );
or2  gate( .a(EX296), .b(EX299), .O(EX300) );
or2  gate( .a(EX298), .b(EX300), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );
inv1 gate( .a(N360),.O(N360_NOT) );
inv1 gate( .a(N27),.O(N27_NOT));
and2 gate( .a(N360_NOT), .b(p121), .O(EX301) );
and2 gate( .a(N27_NOT), .b(EX301), .O(EX302) );
and2 gate( .a(N360), .b(p122), .O(EX303) );
and2 gate( .a(N27_NOT), .b(EX303), .O(EX304) );
and2 gate( .a(N360_NOT), .b(p123), .O(EX305) );
and2 gate( .a(N27), .b(EX305), .O(EX306) );
and2 gate( .a(N360), .b(p124), .O(EX307) );
and2 gate( .a(N27), .b(EX307), .O(EX308) );
or2  gate( .a(EX302), .b(EX304), .O(EX309) );
or2  gate( .a(EX306), .b(EX309), .O(EX310) );
or2  gate( .a(EX308), .b(EX310), .O(N372) );
nand2 gate131( .a(N360), .b(N40), .O(N373) );
nand2 gate132( .a(N360), .b(N53), .O(N374) );
inv1 gate( .a(N360),.O(N360_NOT) );
inv1 gate( .a(N66),.O(N66_NOT));
and2 gate( .a(N360_NOT), .b(p125), .O(EX311) );
and2 gate( .a(N66_NOT), .b(EX311), .O(EX312) );
and2 gate( .a(N360), .b(p126), .O(EX313) );
and2 gate( .a(N66_NOT), .b(EX313), .O(EX314) );
and2 gate( .a(N360_NOT), .b(p127), .O(EX315) );
and2 gate( .a(N66), .b(EX315), .O(EX316) );
and2 gate( .a(N360), .b(p128), .O(EX317) );
and2 gate( .a(N66), .b(EX317), .O(EX318) );
or2  gate( .a(EX312), .b(EX314), .O(EX319) );
or2  gate( .a(EX316), .b(EX319), .O(EX320) );
or2  gate( .a(EX318), .b(EX320), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );
inv1 gate( .a(N360),.O(N360_NOT) );
inv1 gate( .a(N105),.O(N105_NOT));
and2 gate( .a(N360_NOT), .b(p129), .O(EX321) );
and2 gate( .a(N105_NOT), .b(EX321), .O(EX322) );
and2 gate( .a(N360), .b(p130), .O(EX323) );
and2 gate( .a(N105_NOT), .b(EX323), .O(EX324) );
and2 gate( .a(N360_NOT), .b(p131), .O(EX325) );
and2 gate( .a(N105), .b(EX325), .O(EX326) );
and2 gate( .a(N360), .b(p132), .O(EX327) );
and2 gate( .a(N105), .b(EX327), .O(EX328) );
or2  gate( .a(EX322), .b(EX324), .O(EX329) );
or2  gate( .a(EX326), .b(EX329), .O(EX330) );
or2  gate( .a(EX328), .b(EX330), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule
