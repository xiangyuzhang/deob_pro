
module c1908 (N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
              N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
              N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
              N94,N99,N104,N2753,N2754,N2755,N2756,N2762,N2767,N2768,
              N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,
              N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2899);

input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,
      N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
      N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,
      N94,N99,N104;

input p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,
        p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,
        p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,
        p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,
        p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,
        p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,
        p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,
        p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,
        p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,
        p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,
        p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,
        p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,
        p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,
        p131,p132,p133,p134,p135,p136,p137,p138,p139,p140,
        p141,p142,p143,p144,p145,p146,p147,p148,p149,p150,
        p151,p152,p153,p154,p155,p156,p157,p158,p159,p160,
        p161,p162,p163,p164,p165,p166,p167,p168,p169,p170,
        p171,p172,p173,p174,p175,p176,p177,p178,p179,p180,
        p181,p182,p183,p184,p185,p186,p187,p188,p189,p190,
        p191,p192,p193,p194,p195,p196,p197,p198,p199,p200,
        p201,p202,p203,p204,p205,p206,p207,p208,p209,p210,
        p211,p212,p213,p214,p215,p216,p217,p218,p219,p220,
        p221,p222,p223,p224,p225,p226,p227,p228,p229,p230,
        p231,p232,p233,p234,p235,p236,p237,p238,p239,p240,
        p241,p242,p243,p244,p245,p246,p247,p248,p249,p250,
        p251,p252,p253,p254,p255,p256,p257,p258,p259,p260,
        p261,p262,p263,p264,p265,p266,p267,p268,p269,p270,
        p271,p272,p273,p274,p275,p276,p277,p278,p279,p280,
        p281,p282,p283,p284,p285,p286,p287,p288,p289,p290,
        p291,p292,p293,p294,p295,p296,p297,p298,p299,p300,
        p301,p302,p303,p304,p305,p306,p307,p308,p309,p310,
        p311,p312,p313,p314,p315,p316,p317,p318,p319,p320,
        p321,p322,p323,p324,p325,p326,p327,p328,p329,p330,
        p331,p332,p333,p334,p335,p336,p337,p338,p339,p340,
        p341,p342,p343,p344,p345,p346,p347,p348,p349,p350,
        p351,p352,p353,p354,p355,p356,p357,p358,p359,p360,
        p361,p362,p363,p364,p365,p366,p367,p368,p369,p370,
        p371,p372,p373,p374,p375,p376,p377,p378,p379,p380,
        p381,p382,p383,p384,p385,p386,p387,p388,p389,p390,
        p391,p392,p393,p394,p395,p396,p397,p398,p399,p400,
        p401,p402,p403,p404,p405,p406,p407,p408,p409,p410,
        p411,p412,p413,p414,p415,p416,p417,p418,p419,p420;

output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,
       N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
       N2889,N2890,N2891,N2892,N2899;

wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,
     N229,N232,N235,N239,N243,N247,N251,N252,N253,N256,
     N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,
     N283,N290,N297,N300,N303,N306,N313,N316,N319,N326,
     N331,N338,N343,N346,N349,N352,N355,N358,N361,N364,
     N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,
     N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
     N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
     N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,
     N586,N589,N592,N595,N598,N601,N602,N603,N608,N612,
     N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,
     N646,N649,N652,N655,N658,N661,N664,N667,N670,N673,
     N676,N679,N682,N685,N688,N691,N694,N697,N700,N703,
     N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,
     N736,N739,N742,N745,N748,N751,N886,N887,N888,N889,
     N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
     N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,
     N920,N921,N922,N923,N926,N935,N938,N939,N942,N943,
     N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,
     N968,N969,N972,N973,N976,N977,N980,N981,N984,N985,
     N988,N989,N990,N991,N992,N993,N994,N997,N998,N1001,
     N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,
     N1016,N1019,N1022,N1025,N1028,N1031,N1034,N1037,N1040,N1043,
     N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
     N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,
     N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,
     N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,
     N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
     N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,
     N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,
     N1240,N1241,N1242,N1243,N1246,N1249,N1252,N1255,N1258,N1261,
     N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
     N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,
     N1348,N1349,N1350,N1351,N1352,N1355,N1358,N1361,N1364,N1367,
     N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,
     N1393,N1396,N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,
     N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447,
     N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,
     N1460,N1461,N1462,N1463,N1464,N1468,N1469,N1470,N1471,N1472,
     N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
     N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,
     N1510,N1513,N1514,N1517,N1520,N1521,N1522,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,
     N1561,N1567,N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,
     N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,N1620,N1623,
     N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,
     N1664,N1671,N1672,N1675,N1677,N1678,N1679,N1680,N1681,N1682,
     N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
     N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,
     N1730,N1731,N1734,N1740,N1741,N1742,N1746,N1747,N1748,N1751,
     N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,
     N1777,N1783,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,
     N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,N1812,N1815,
     N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,
     N1838,N1841,N1848,N1849,N1850,N1852,N1855,N1856,N1857,N1858,
     N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
     N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,
     N1912,N1913,N1915,N1919,N1920,N1921,N1922,N1923,N1924,N1927,
     N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,
     N1953,N1958,N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,
     N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,N2005,N2006,
     N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,
     N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2030,N2033,
     N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
     N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,
     N2086,N2089,N2104,N2119,N2129,N2143,N2148,N2151,N2196,N2199,
     N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,
     N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
     N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,N2256,N2257,
     N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,
     N2340,N2353,N2361,N2375,N2384,N2385,N2386,N2426,N2427,N2537,
     N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
     N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,
     N2617,N2620,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,
     N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,
     N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,
     N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,N2724,N2725,
     N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,
     N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,
     N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
     N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,
     N2810,N2812,N2815,N2818,N2821,N2824,N2827,N2828,N2829,N2843,
     N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,
     N2861,N2862,N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
     N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,
     N2883,N2895,N2896,N2897,N2898,
     N66_NOT,N91_NOT,N306_NOT,N331_NOT,N306_NOT,N331_NOT,N306_NOT,N331_NOT,N63_NOT,N319_NOT,
     N260_NOT,N72_NOT,N256_NOT,N300_NOT,N252_NOT,N316_NOT,N56_NOT,N608_NOT,N616_NOT,N889_NOT,
     N622_NOT,N891_NOT,N655_NOT,N895_NOT,N652_NOT,N896_NOT,N727_NOT,N991_NOT,N739_NOT,N1002_NOT,
     N748_NOT,N1009_NOT,N1054_NOT,N1055_NOT,N985_NOT,N892_NOT,N922_NOT,N923_NOT,N981_NOT,N984_NOT,
     N1049_NOT,N1001_NOT,N1132_NOT,N1133_NOT,N709_NOT,N1223_NOT,N712_NOT,N1225_NOT,N628_NOT,N1230_NOT,
     N730_NOT,N1238_NOT,N1267_NOT,N1160_NOT,N1311_NOT,N1210_NOT,N1312_NOT,N1212_NOT,N1317_NOT,N1226_NOT,
     N1322_NOT,N1231_NOT,N1232_NOT,N990_NOT,N1235_NOT,N993_NOT,N649_NOT,N1346_NOT,N637_NOT,N1388_NOT,
     N1352_NOT,N1149_NOT,N1361_NOT,N1152_NOT,N1379_NOT,N1157_NOT,N1376_NOT,N1227_NOT,N1397_NOT,N1438_NOT,
     N939_NOT,N1444_NOT,N935_NOT,N1446_NOT,N998_NOT,N1463_NOT,N965_NOT,N1468_NOT,N1453_NOT,N1493_NOT,
     N1455_NOT,N1494_NOT,N1476_NOT,N1504_NOT,N1481_NOT,N1532_NOT,N1567_NOT,N1568_NOT,N1478_NOT,N1595_NOT,
     N1594_NOT,N1636_NOT,N1510_NOT,N1639_NOT,N1647_NOT,N1675_NOT,N1031_NOT,N1681_NOT,N1658_NOT,N1593_NOT,
     N1638_NOT,N1688_NOT,N1685_NOT,N1528_NOT,N1600_NOT,N1709_NOT,N1678_NOT,N1712_NOT,N1537_NOT,N1721_NOT,
     N1697_NOT,N1727_NOT,N1708_NOT,N1746_NOT,N1664_NOT,N1763_NOT,N1334_NOT,N1773_NOT,N1777_NOT,N1490_NOT,
     N1815_NOT,N1707_NOT,N1855_NOT,N1885_NOT,N679_NOT,N1920_NOT,N676_NOT,N1922_NOT,N1921_NOT,N1942_NOT,
     N1947_NOT,N1499_NOT,N673_NOT,N1976_NOT,N1258_NOT,N2007_NOT,N1977_NOT,N2009_NOT,N1534_NOT,N2021_NOT,
     N2004_NOT,N2024_NOT,N2060_NOT,N290_NOT,N2199_NOT,N1348_NOT,N2196_NOT,N1349_NOT,N667_NOT,N2215_NOT,
     N664_NOT,N2217_NOT,N1255_NOT,N2223_NOT,N1252_NOT,N2225_NOT,N2228_NOT,N2235_NOT,N1164_NOT,N2241_NOT,
     N1168_NOT,N2245_NOT,N2089_NOT,N2260_NOT,N1164_NOT,N2263_NOT,N2567_NOT,N537_NOT,N352_NOT,N2676_NOT,
     N370_NOT,N2683_NOT,N2673_NOT,N2722_NOT,N361_NOT,N2729_NOT,N364_NOT,N2731_NOT,N379_NOT,N2740_NOT,
     N2776_NOT,N2019_NOT,N2384_NOT,N2800_NOT,N2829_NOT,N1985_NOT,N1866_NOT,N2859_NOT,N1902_NOT,N2861_NOT,
     N2843_NOT,N886_NOT,N2846_NOT,N887_NOT,N685_NOT,N2874_NOT,N2871_NOT,N2881_NOT,N2895_NOT,N2897_NOT,
     EX1,EX2,EX3,EX4,EX5,EX6,EX7,EX8,EX9,EX10,
     EX11,EX12,EX13,EX14,EX15,EX16,EX17,EX18,EX19,EX20,
     EX21,EX22,EX23,EX24,EX25,EX26,EX27,EX28,EX29,EX30,
     EX31,EX32,EX33,EX34,EX35,EX36,EX37,EX38,EX39,EX40,
     EX41,EX42,EX43,EX44,EX45,EX46,EX47,EX48,EX49,EX50,
     EX51,EX52,EX53,EX54,EX55,EX56,EX57,EX58,EX59,EX60,
     EX61,EX62,EX63,EX64,EX65,EX66,EX67,EX68,EX69,EX70,
     EX71,EX72,EX73,EX74,EX75,EX76,EX77,EX78,EX79,EX80,
     EX81,EX82,EX83,EX84,EX85,EX86,EX87,EX88,EX89,EX90,
     EX91,EX92,EX93,EX94,EX95,EX96,EX97,EX98,EX99,EX100,
     EX101,EX102,EX103,EX104,EX105,EX106,EX107,EX108,EX109,EX110,
     EX111,EX112,EX113,EX114,EX115,EX116,EX117,EX118,EX119,EX120,
     EX121,EX122,EX123,EX124,EX125,EX126,EX127,EX128,EX129,EX130,
     EX131,EX132,EX133,EX134,EX135,EX136,EX137,EX138,EX139,EX140,
     EX141,EX142,EX143,EX144,EX145,EX146,EX147,EX148,EX149,EX150,
     EX151,EX152,EX153,EX154,EX155,EX156,EX157,EX158,EX159,EX160,
     EX161,EX162,EX163,EX164,EX165,EX166,EX167,EX168,EX169,EX170,
     EX171,EX172,EX173,EX174,EX175,EX176,EX177,EX178,EX179,EX180,
     EX181,EX182,EX183,EX184,EX185,EX186,EX187,EX188,EX189,EX190,
     EX191,EX192,EX193,EX194,EX195,EX196,EX197,EX198,EX199,EX200,
     EX201,EX202,EX203,EX204,EX205,EX206,EX207,EX208,EX209,EX210,
     EX211,EX212,EX213,EX214,EX215,EX216,EX217,EX218,EX219,EX220,
     EX221,EX222,EX223,EX224,EX225,EX226,EX227,EX228,EX229,EX230,
     EX231,EX232,EX233,EX234,EX235,EX236,EX237,EX238,EX239,EX240,
     EX241,EX242,EX243,EX244,EX245,EX246,EX247,EX248,EX249,EX250,
     EX251,EX252,EX253,EX254,EX255,EX256,EX257,EX258,EX259,EX260,
     EX261,EX262,EX263,EX264,EX265,EX266,EX267,EX268,EX269,EX270,
     EX271,EX272,EX273,EX274,EX275,EX276,EX277,EX278,EX279,EX280,
     EX281,EX282,EX283,EX284,EX285,EX286,EX287,EX288,EX289,EX290,
     EX291,EX292,EX293,EX294,EX295,EX296,EX297,EX298,EX299,EX300,
     EX301,EX302,EX303,EX304,EX305,EX306,EX307,EX308,EX309,EX310,
     EX311,EX312,EX313,EX314,EX315,EX316,EX317,EX318,EX319,EX320,
     EX321,EX322,EX323,EX324,EX325,EX326,EX327,EX328,EX329,EX330,
     EX331,EX332,EX333,EX334,EX335,EX336,EX337,EX338,EX339,EX340,
     EX341,EX342,EX343,EX344,EX345,EX346,EX347,EX348,EX349,EX350,
     EX351,EX352,EX353,EX354,EX355,EX356,EX357,EX358,EX359,EX360,
     EX361,EX362,EX363,EX364,EX365,EX366,EX367,EX368,EX369,EX370,
     EX371,EX372,EX373,EX374,EX375,EX376,EX377,EX378,EX379,EX380,
     EX381,EX382,EX383,EX384,EX385,EX386,EX387,EX388,EX389,EX390,
     EX391,EX392,EX393,EX394,EX395,EX396,EX397,EX398,EX399,EX400,
     EX401,EX402,EX403,EX404,EX405,EX406,EX407,EX408,EX409,EX410,
     EX411,EX412,EX413,EX414,EX415,EX416,EX417,EX418,EX419,EX420,
     EX421,EX422,EX423,EX424,EX425,EX426,EX427,EX428,EX429,EX430,
     EX431,EX432,EX433,EX434,EX435,EX436,EX437,EX438,EX439,EX440,
     EX441,EX442,EX443,EX444,EX445,EX446,EX447,EX448,EX449,EX450,
     EX451,EX452,EX453,EX454,EX455,EX456,EX457,EX458,EX459,EX460,
     EX461,EX462,EX463,EX464,EX465,EX466,EX467,EX468,EX469,EX470,
     EX471,EX472,EX473,EX474,EX475,EX476,EX477,EX478,EX479,EX480,
     EX481,EX482,EX483,EX484,EX485,EX486,EX487,EX488,EX489,EX490,
     EX491,EX492,EX493,EX494,EX495,EX496,EX497,EX498,EX499,EX500,
     EX501,EX502,EX503,EX504,EX505,EX506,EX507,EX508,EX509,EX510,
     EX511,EX512,EX513,EX514,EX515,EX516,EX517,EX518,EX519,EX520,
     EX521,EX522,EX523,EX524,EX525,EX526,EX527,EX528,EX529,EX530,
     EX531,EX532,EX533,EX534,EX535,EX536,EX537,EX538,EX539,EX540,
     EX541,EX542,EX543,EX544,EX545,EX546,EX547,EX548,EX549,EX550,
     EX551,EX552,EX553,EX554,EX555,EX556,EX557,EX558,EX559,EX560,
     EX561,EX562,EX563,EX564,EX565,EX566,EX567,EX568,EX569,EX570,
     EX571,EX572,EX573,EX574,EX575,EX576,EX577,EX578,EX579,EX580,
     EX581,EX582,EX583,EX584,EX585,EX586,EX587,EX588,EX589,EX590,
     EX591,EX592,EX593,EX594,EX595,EX596,EX597,EX598,EX599,EX600,
     EX601,EX602,EX603,EX604,EX605,EX606,EX607,EX608,EX609,EX610,
     EX611,EX612,EX613,EX614,EX615,EX616,EX617,EX618,EX619,EX620,
     EX621,EX622,EX623,EX624,EX625,EX626,EX627,EX628,EX629,EX630,
     EX631,EX632,EX633,EX634,EX635,EX636,EX637,EX638,EX639,EX640,
     EX641,EX642,EX643,EX644,EX645,EX646,EX647,EX648,EX649,EX650,
     EX651,EX652,EX653,EX654,EX655,EX656,EX657,EX658,EX659,EX660,
     EX661,EX662,EX663,EX664,EX665,EX666,EX667,EX668,EX669,EX670,
     EX671,EX672,EX673,EX674,EX675,EX676,EX677,EX678,EX679,EX680,
     EX681,EX682,EX683,EX684,EX685,EX686,EX687,EX688,EX689,EX690,
     EX691,EX692,EX693,EX694,EX695,EX696,EX697,EX698,EX699,EX700,
     EX701,EX702,EX703,EX704,EX705,EX706,EX707,EX708,EX709,EX710,
     EX711,EX712,EX713,EX714,EX715,EX716,EX717,EX718,EX719,EX720,
     EX721,EX722,EX723,EX724,EX725,EX726,EX727,EX728,EX729,EX730,
     EX731,EX732,EX733,EX734,EX735,EX736,EX737,EX738,EX739,EX740,
     EX741,EX742,EX743,EX744,EX745,EX746,EX747,EX748,EX749,EX750,
     EX751,EX752,EX753,EX754,EX755,EX756,EX757,EX758,EX759,EX760,
     EX761,EX762,EX763,EX764,EX765,EX766,EX767,EX768,EX769,EX770,
     EX771,EX772,EX773,EX774,EX775,EX776,EX777,EX778,EX779,EX780,
     EX781,EX782,EX783,EX784,EX785,EX786,EX787,EX788,EX789,EX790,
     EX791,EX792,EX793,EX794,EX795,EX796,EX797,EX798,EX799,EX800,
     EX801,EX802,EX803,EX804,EX805,EX806,EX807,EX808,EX809,EX810,
     EX811,EX812,EX813,EX814,EX815,EX816,EX817,EX818,EX819,EX820,
     EX821,EX822,EX823,EX824,EX825,EX826,EX827,EX828,EX829,EX830,
     EX831,EX832,EX833,EX834,EX835,EX836,EX837,EX838,EX839,EX840,
     EX841,EX842,EX843,EX844,EX845,EX846,EX847,EX848,EX849,EX850,
     EX851,EX852,EX853,EX854,EX855,EX856,EX857,EX858,EX859,EX860,
     EX861,EX862,EX863,EX864,EX865,EX866,EX867,EX868,EX869,EX870,
     EX871,EX872,EX873,EX874,EX875,EX876,EX877,EX878,EX879,EX880,
     EX881,EX882,EX883,EX884,EX885,EX886,EX887,EX888,EX889,EX890,
     EX891,EX892,EX893,EX894,EX895,EX896,EX897,EX898,EX899,EX900,
     EX901,EX902,EX903,EX904,EX905,EX906,EX907,EX908,EX909,EX910,
     EX911,EX912,EX913,EX914,EX915,EX916,EX917,EX918,EX919,EX920,
     EX921,EX922,EX923,EX924,EX925,EX926,EX927,EX928,EX929,EX930,
     EX931,EX932,EX933,EX934,EX935,EX936,EX937,EX938,EX939,EX940,
     EX941,EX942,EX943,EX944,EX945,EX946,EX947,EX948,EX949,EX950,
     EX951,EX952,EX953,EX954,EX955,EX956,EX957,EX958,EX959,EX960,
     EX961,EX962,EX963,EX964,EX965,EX966,EX967,EX968,EX969,EX970,
     EX971,EX972,EX973,EX974,EX975,EX976,EX977,EX978,EX979,EX980,
     EX981,EX982,EX983,EX984,EX985,EX986,EX987,EX988,EX989,EX990,
     EX991,EX992,EX993,EX994,EX995,EX996,EX997,EX998,EX999,EX1000,
     EX1001,EX1002,EX1003,EX1004,EX1005,EX1006,EX1007,EX1008,EX1009,EX1010,
     EX1011,EX1012,EX1013,EX1014,EX1015,EX1016,EX1017,EX1018,EX1019,EX1020,
     EX1021,EX1022,EX1023,EX1024,EX1025,EX1026,EX1027,EX1028,EX1029,EX1030,
     EX1031,EX1032,EX1033,EX1034,EX1035,EX1036,EX1037,EX1038,EX1039,EX1040,
     EX1041,EX1042,EX1043,EX1044,EX1045,EX1046,EX1047,EX1048,EX1049,EX1050;


inv1 gate1( .a(N1), .O(N190) );
inv1 gate2( .a(N4), .O(N194) );
inv1 gate3( .a(N7), .O(N197) );
inv1 gate4( .a(N10), .O(N201) );
inv1 gate5( .a(N13), .O(N206) );
inv1 gate6( .a(N16), .O(N209) );
inv1 gate7( .a(N19), .O(N212) );
inv1 gate8( .a(N22), .O(N216) );
inv1 gate9( .a(N25), .O(N220) );
inv1 gate10( .a(N28), .O(N225) );
inv1 gate11( .a(N31), .O(N229) );
inv1 gate12( .a(N34), .O(N232) );
inv1 gate13( .a(N37), .O(N235) );
inv1 gate14( .a(N40), .O(N239) );
inv1 gate15( .a(N43), .O(N243) );
inv1 gate16( .a(N46), .O(N247) );
nand2 gate17( .a(N63), .b(N88), .O(N251) );
inv1 gate( .a(N66),.O(N66_NOT) );
inv1 gate( .a(N91),.O(N91_NOT));
and2 gate( .a(N66_NOT), .b(p1), .O(EX1) );
and2 gate( .a(N91_NOT), .b(EX1), .O(EX2) );
and2 gate( .a(N66), .b(p2), .O(EX3) );
and2 gate( .a(N91_NOT), .b(EX3), .O(EX4) );
and2 gate( .a(N66_NOT), .b(p3), .O(EX5) );
and2 gate( .a(N91), .b(EX5), .O(EX6) );
and2 gate( .a(N66), .b(p4), .O(EX7) );
and2 gate( .a(N91), .b(EX7), .O(EX8) );
or2  gate( .a(EX2), .b(EX4), .O(EX9) );
or2  gate( .a(EX6), .b(EX9), .O(EX10) );
or2  gate( .a(EX8), .b(EX10), .O(N252) );
inv1 gate19( .a(N72), .O(N253) );
inv1 gate20( .a(N72), .O(N256) );
buf1 gate21( .a(N69), .O(N257) );
buf1 gate22( .a(N69), .O(N260) );
inv1 gate23( .a(N76), .O(N263) );
inv1 gate24( .a(N79), .O(N266) );
inv1 gate25( .a(N82), .O(N269) );
inv1 gate26( .a(N85), .O(N272) );
inv1 gate27( .a(N104), .O(N275) );
inv1 gate28( .a(N104), .O(N276) );
inv1 gate29( .a(N88), .O(N277) );
inv1 gate30( .a(N91), .O(N280) );
buf1 gate31( .a(N94), .O(N283) );
inv1 gate32( .a(N94), .O(N290) );
buf1 gate33( .a(N94), .O(N297) );
inv1 gate34( .a(N94), .O(N300) );
buf1 gate35( .a(N99), .O(N303) );
inv1 gate36( .a(N99), .O(N306) );
inv1 gate37( .a(N99), .O(N313) );
buf1 gate38( .a(N104), .O(N316) );
inv1 gate39( .a(N104), .O(N319) );
buf1 gate40( .a(N104), .O(N326) );
buf1 gate41( .a(N104), .O(N331) );
inv1 gate42( .a(N104), .O(N338) );
buf1 gate43( .a(N1), .O(N343) );
buf1 gate44( .a(N4), .O(N346) );
buf1 gate45( .a(N7), .O(N349) );
buf1 gate46( .a(N10), .O(N352) );
buf1 gate47( .a(N13), .O(N355) );
buf1 gate48( .a(N16), .O(N358) );
buf1 gate49( .a(N19), .O(N361) );
buf1 gate50( .a(N22), .O(N364) );
buf1 gate51( .a(N25), .O(N367) );
buf1 gate52( .a(N28), .O(N370) );
buf1 gate53( .a(N31), .O(N373) );
buf1 gate54( .a(N34), .O(N376) );
buf1 gate55( .a(N37), .O(N379) );
buf1 gate56( .a(N40), .O(N382) );
buf1 gate57( .a(N43), .O(N385) );
buf1 gate58( .a(N46), .O(N388) );
inv1 gate59( .a(N343), .O(N534) );
inv1 gate60( .a(N346), .O(N535) );
inv1 gate61( .a(N349), .O(N536) );
inv1 gate62( .a(N352), .O(N537) );
inv1 gate63( .a(N355), .O(N538) );
inv1 gate64( .a(N358), .O(N539) );
inv1 gate65( .a(N361), .O(N540) );
inv1 gate66( .a(N364), .O(N541) );
inv1 gate67( .a(N367), .O(N542) );
inv1 gate68( .a(N370), .O(N543) );
inv1 gate69( .a(N373), .O(N544) );
inv1 gate70( .a(N376), .O(N545) );
inv1 gate71( .a(N379), .O(N546) );
inv1 gate72( .a(N382), .O(N547) );
inv1 gate73( .a(N385), .O(N548) );
inv1 gate74( .a(N388), .O(N549) );
inv1 gate( .a(N306),.O(N306_NOT) );
inv1 gate( .a(N331),.O(N331_NOT));
and2 gate( .a(N306_NOT), .b(p5), .O(EX11) );
and2 gate( .a(N331_NOT), .b(EX11), .O(EX12) );
and2 gate( .a(N306), .b(p6), .O(EX13) );
and2 gate( .a(N331_NOT), .b(EX13), .O(EX14) );
and2 gate( .a(N306_NOT), .b(p7), .O(EX15) );
and2 gate( .a(N331), .b(EX15), .O(EX16) );
and2 gate( .a(N306), .b(p8), .O(EX17) );
and2 gate( .a(N331), .b(EX17), .O(EX18) );
or2  gate( .a(EX12), .b(EX14), .O(EX19) );
or2  gate( .a(EX16), .b(EX19), .O(EX20) );
or2  gate( .a(EX18), .b(EX20), .O(N550) );
nand2 gate76( .a(N306), .b(N331), .O(N551) );
nand2 gate77( .a(N306), .b(N331), .O(N552) );
inv1 gate( .a(N306),.O(N306_NOT) );
inv1 gate( .a(N331),.O(N331_NOT));
and2 gate( .a(N306_NOT), .b(p9), .O(EX21) );
and2 gate( .a(N331_NOT), .b(EX21), .O(EX22) );
and2 gate( .a(N306), .b(p10), .O(EX23) );
and2 gate( .a(N331_NOT), .b(EX23), .O(EX24) );
and2 gate( .a(N306_NOT), .b(p11), .O(EX25) );
and2 gate( .a(N331), .b(EX25), .O(EX26) );
and2 gate( .a(N306), .b(p12), .O(EX27) );
and2 gate( .a(N331), .b(EX27), .O(EX28) );
or2  gate( .a(EX22), .b(EX24), .O(EX29) );
or2  gate( .a(EX26), .b(EX29), .O(EX30) );
or2  gate( .a(EX28), .b(EX30), .O(N553) );
nand2 gate79( .a(N306), .b(N331), .O(N554) );
inv1 gate( .a(N306),.O(N306_NOT) );
inv1 gate( .a(N331),.O(N331_NOT));
and2 gate( .a(N306_NOT), .b(p13), .O(EX31) );
and2 gate( .a(N331_NOT), .b(EX31), .O(EX32) );
and2 gate( .a(N306), .b(p14), .O(EX33) );
and2 gate( .a(N331_NOT), .b(EX33), .O(EX34) );
and2 gate( .a(N306_NOT), .b(p15), .O(EX35) );
and2 gate( .a(N331), .b(EX35), .O(EX36) );
and2 gate( .a(N306), .b(p16), .O(EX37) );
and2 gate( .a(N331), .b(EX37), .O(EX38) );
or2  gate( .a(EX32), .b(EX34), .O(EX39) );
or2  gate( .a(EX36), .b(EX39), .O(EX40) );
or2  gate( .a(EX38), .b(EX40), .O(N555) );
buf1 gate81( .a(N190), .O(N556) );
buf1 gate82( .a(N194), .O(N559) );
buf1 gate83( .a(N206), .O(N562) );
buf1 gate84( .a(N209), .O(N565) );
buf1 gate85( .a(N225), .O(N568) );
buf1 gate86( .a(N243), .O(N571) );
inv1 gate( .a(N63),.O(N63_NOT) );
inv1 gate( .a(N319),.O(N319_NOT));
and2 gate( .a(N63_NOT), .b(p17), .O(EX41) );
and2 gate( .a(N319_NOT), .b(EX41), .O(EX42) );
and2 gate( .a(N63), .b(p18), .O(EX43) );
and2 gate( .a(N319_NOT), .b(EX43), .O(EX44) );
and2 gate( .a(N63_NOT), .b(p19), .O(EX45) );
and2 gate( .a(N319), .b(EX45), .O(EX46) );
and2 gate( .a(N63), .b(p20), .O(EX47) );
and2 gate( .a(N319), .b(EX47), .O(EX48) );
or2  gate( .a(EX42), .b(EX44), .O(EX49) );
or2  gate( .a(EX46), .b(EX49), .O(EX50) );
or2  gate( .a(EX48), .b(EX50), .O(N574) );
buf1 gate88( .a(N220), .O(N577) );
buf1 gate89( .a(N229), .O(N580) );
buf1 gate90( .a(N232), .O(N583) );
and2 gate91( .a(N66), .b(N319), .O(N586) );
buf1 gate92( .a(N239), .O(N589) );
and3 gate93( .a(N49), .b(N253), .c(N319), .O(N592) );
buf1 gate94( .a(N247), .O(N595) );
buf1 gate95( .a(N239), .O(N598) );
nand2 gate96( .a(N326), .b(N277), .O(N601) );
nand2 gate97( .a(N326), .b(N280), .O(N602) );
inv1 gate( .a(N260),.O(N260_NOT) );
inv1 gate( .a(N72),.O(N72_NOT));
and2 gate( .a(N260_NOT), .b(p21), .O(EX51) );
and2 gate( .a(N72_NOT), .b(EX51), .O(EX52) );
and2 gate( .a(N260), .b(p22), .O(EX53) );
and2 gate( .a(N72_NOT), .b(EX53), .O(EX54) );
and2 gate( .a(N260_NOT), .b(p23), .O(EX55) );
and2 gate( .a(N72), .b(EX55), .O(EX56) );
and2 gate( .a(N260), .b(p24), .O(EX57) );
and2 gate( .a(N72), .b(EX57), .O(EX58) );
or2  gate( .a(EX52), .b(EX54), .O(EX59) );
or2  gate( .a(EX56), .b(EX59), .O(EX60) );
or2  gate( .a(EX58), .b(EX60), .O(N603) );
nand2 gate99( .a(N260), .b(N300), .O(N608) );
inv1 gate( .a(N256),.O(N256_NOT) );
inv1 gate( .a(N300),.O(N300_NOT));
and2 gate( .a(N256_NOT), .b(p25), .O(EX61) );
and2 gate( .a(N300_NOT), .b(EX61), .O(EX62) );
and2 gate( .a(N256), .b(p26), .O(EX63) );
and2 gate( .a(N300_NOT), .b(EX63), .O(EX64) );
and2 gate( .a(N256_NOT), .b(p27), .O(EX65) );
and2 gate( .a(N300), .b(EX65), .O(EX66) );
and2 gate( .a(N256), .b(p28), .O(EX67) );
and2 gate( .a(N300), .b(EX67), .O(EX68) );
or2  gate( .a(EX62), .b(EX64), .O(EX69) );
or2  gate( .a(EX66), .b(EX69), .O(EX70) );
or2  gate( .a(EX68), .b(EX70), .O(N612) );
buf1 gate101( .a(N201), .O(N616) );
buf1 gate102( .a(N216), .O(N619) );
buf1 gate103( .a(N220), .O(N622) );
buf1 gate104( .a(N239), .O(N625) );
buf1 gate105( .a(N190), .O(N628) );
buf1 gate106( .a(N190), .O(N631) );
buf1 gate107( .a(N194), .O(N634) );
buf1 gate108( .a(N229), .O(N637) );
buf1 gate109( .a(N197), .O(N640) );
and3 gate110( .a(N56), .b(N257), .c(N319), .O(N643) );
buf1 gate111( .a(N232), .O(N646) );
buf1 gate112( .a(N201), .O(N649) );
buf1 gate113( .a(N235), .O(N652) );
and3 gate114( .a(N60), .b(N257), .c(N319), .O(N655) );
buf1 gate115( .a(N263), .O(N658) );
buf1 gate116( .a(N263), .O(N661) );
buf1 gate117( .a(N266), .O(N664) );
buf1 gate118( .a(N266), .O(N667) );
buf1 gate119( .a(N269), .O(N670) );
buf1 gate120( .a(N269), .O(N673) );
buf1 gate121( .a(N272), .O(N676) );
buf1 gate122( .a(N272), .O(N679) );
and2 gate123( .a(N251), .b(N316), .O(N682) );
inv1 gate( .a(N252),.O(N252_NOT) );
inv1 gate( .a(N316),.O(N316_NOT));
and2 gate( .a(N252_NOT), .b(p29), .O(EX71) );
and2 gate( .a(N316_NOT), .b(EX71), .O(EX72) );
and2 gate( .a(N252), .b(p30), .O(EX73) );
and2 gate( .a(N316_NOT), .b(EX73), .O(EX74) );
and2 gate( .a(N252_NOT), .b(p31), .O(EX75) );
and2 gate( .a(N316), .b(EX75), .O(EX76) );
and2 gate( .a(N252), .b(p32), .O(EX77) );
and2 gate( .a(N316), .b(EX77), .O(EX78) );
or2  gate( .a(EX72), .b(EX74), .O(EX79) );
or2  gate( .a(EX76), .b(EX79), .O(EX80) );
or2  gate( .a(EX78), .b(EX80), .O(N685) );
buf1 gate125( .a(N197), .O(N688) );
buf1 gate126( .a(N197), .O(N691) );
buf1 gate127( .a(N212), .O(N694) );
buf1 gate128( .a(N212), .O(N697) );
buf1 gate129( .a(N247), .O(N700) );
buf1 gate130( .a(N247), .O(N703) );
buf1 gate131( .a(N235), .O(N706) );
buf1 gate132( .a(N235), .O(N709) );
buf1 gate133( .a(N201), .O(N712) );
buf1 gate134( .a(N201), .O(N715) );
buf1 gate135( .a(N206), .O(N718) );
buf1 gate136( .a(N216), .O(N721) );
and3 gate137( .a(N53), .b(N253), .c(N319), .O(N724) );
buf1 gate138( .a(N243), .O(N727) );
buf1 gate139( .a(N220), .O(N730) );
buf1 gate140( .a(N220), .O(N733) );
buf1 gate141( .a(N209), .O(N736) );
buf1 gate142( .a(N216), .O(N739) );
buf1 gate143( .a(N225), .O(N742) );
buf1 gate144( .a(N243), .O(N745) );
buf1 gate145( .a(N212), .O(N748) );
buf1 gate146( .a(N225), .O(N751) );
inv1 gate147( .a(N682), .O(N886) );
inv1 gate148( .a(N685), .O(N887) );
inv1 gate149( .a(N616), .O(N888) );
inv1 gate150( .a(N619), .O(N889) );
inv1 gate151( .a(N622), .O(N890) );
inv1 gate152( .a(N625), .O(N891) );
inv1 gate153( .a(N631), .O(N892) );
inv1 gate154( .a(N643), .O(N893) );
inv1 gate155( .a(N649), .O(N894) );
inv1 gate156( .a(N652), .O(N895) );
inv1 gate157( .a(N655), .O(N896) );
and2 gate158( .a(N49), .b(N612), .O(N897) );
and2 gate159( .a(N56), .b(N608), .O(N898) );
nand2 gate160( .a(N53), .b(N612), .O(N899) );
nand2 gate161( .a(N60), .b(N608), .O(N903) );
nand2 gate162( .a(N49), .b(N612), .O(N907) );
inv1 gate( .a(N56),.O(N56_NOT) );
inv1 gate( .a(N608),.O(N608_NOT));
and2 gate( .a(N56_NOT), .b(p33), .O(EX81) );
and2 gate( .a(N608_NOT), .b(EX81), .O(EX82) );
and2 gate( .a(N56), .b(p34), .O(EX83) );
and2 gate( .a(N608_NOT), .b(EX83), .O(EX84) );
and2 gate( .a(N56_NOT), .b(p35), .O(EX85) );
and2 gate( .a(N608), .b(EX85), .O(EX86) );
and2 gate( .a(N56), .b(p36), .O(EX87) );
and2 gate( .a(N608), .b(EX87), .O(EX88) );
or2  gate( .a(EX82), .b(EX84), .O(EX89) );
or2  gate( .a(EX86), .b(EX89), .O(EX90) );
or2  gate( .a(EX88), .b(EX90), .O(N910) );
inv1 gate164( .a(N661), .O(N913) );
inv1 gate165( .a(N658), .O(N914) );
inv1 gate166( .a(N667), .O(N915) );
inv1 gate167( .a(N664), .O(N916) );
inv1 gate168( .a(N673), .O(N917) );
inv1 gate169( .a(N670), .O(N918) );
inv1 gate170( .a(N679), .O(N919) );
inv1 gate171( .a(N676), .O(N920) );
nand4 gate172( .a(N277), .b(N297), .c(N326), .d(N603), .O(N921) );
nand4 gate173( .a(N280), .b(N297), .c(N326), .d(N603), .O(N922) );
nand3 gate174( .a(N303), .b(N338), .c(N603), .O(N923) );
and3 gate175( .a(N303), .b(N338), .c(N603), .O(N926) );
buf1 gate176( .a(N556), .O(N935) );
inv1 gate177( .a(N688), .O(N938) );
buf1 gate178( .a(N556), .O(N939) );
inv1 gate179( .a(N691), .O(N942) );
buf1 gate180( .a(N562), .O(N943) );
inv1 gate181( .a(N694), .O(N946) );
buf1 gate182( .a(N562), .O(N947) );
inv1 gate183( .a(N697), .O(N950) );
buf1 gate184( .a(N568), .O(N951) );
inv1 gate185( .a(N700), .O(N954) );
buf1 gate186( .a(N568), .O(N955) );
inv1 gate187( .a(N703), .O(N958) );
buf1 gate188( .a(N574), .O(N959) );
buf1 gate189( .a(N574), .O(N962) );
buf1 gate190( .a(N580), .O(N965) );
inv1 gate191( .a(N706), .O(N968) );
buf1 gate192( .a(N580), .O(N969) );
inv1 gate193( .a(N709), .O(N972) );
buf1 gate194( .a(N586), .O(N973) );
inv1 gate195( .a(N712), .O(N976) );
buf1 gate196( .a(N586), .O(N977) );
inv1 gate197( .a(N715), .O(N980) );
buf1 gate198( .a(N592), .O(N981) );
inv1 gate199( .a(N628), .O(N984) );
buf1 gate200( .a(N592), .O(N985) );
inv1 gate201( .a(N718), .O(N988) );
inv1 gate202( .a(N721), .O(N989) );
inv1 gate203( .a(N634), .O(N990) );
inv1 gate204( .a(N724), .O(N991) );
inv1 gate205( .a(N727), .O(N992) );
inv1 gate206( .a(N637), .O(N993) );
buf1 gate207( .a(N595), .O(N994) );
inv1 gate208( .a(N730), .O(N997) );
buf1 gate209( .a(N595), .O(N998) );
inv1 gate210( .a(N733), .O(N1001) );
inv1 gate211( .a(N736), .O(N1002) );
inv1 gate212( .a(N739), .O(N1003) );
inv1 gate213( .a(N640), .O(N1004) );
inv1 gate214( .a(N742), .O(N1005) );
inv1 gate215( .a(N745), .O(N1006) );
inv1 gate216( .a(N646), .O(N1007) );
inv1 gate217( .a(N748), .O(N1008) );
inv1 gate218( .a(N751), .O(N1009) );
buf1 gate219( .a(N559), .O(N1010) );
buf1 gate220( .a(N559), .O(N1013) );
buf1 gate221( .a(N565), .O(N1016) );
buf1 gate222( .a(N565), .O(N1019) );
buf1 gate223( .a(N571), .O(N1022) );
buf1 gate224( .a(N571), .O(N1025) );
buf1 gate225( .a(N577), .O(N1028) );
buf1 gate226( .a(N577), .O(N1031) );
buf1 gate227( .a(N583), .O(N1034) );
buf1 gate228( .a(N583), .O(N1037) );
buf1 gate229( .a(N589), .O(N1040) );
buf1 gate230( .a(N589), .O(N1043) );
buf1 gate231( .a(N598), .O(N1046) );
buf1 gate232( .a(N598), .O(N1049) );
nand2 gate233( .a(N619), .b(N888), .O(N1054) );
inv1 gate( .a(N616),.O(N616_NOT) );
inv1 gate( .a(N889),.O(N889_NOT));
and2 gate( .a(N616_NOT), .b(p37), .O(EX91) );
and2 gate( .a(N889_NOT), .b(EX91), .O(EX92) );
and2 gate( .a(N616), .b(p38), .O(EX93) );
and2 gate( .a(N889_NOT), .b(EX93), .O(EX94) );
and2 gate( .a(N616_NOT), .b(p39), .O(EX95) );
and2 gate( .a(N889), .b(EX95), .O(EX96) );
and2 gate( .a(N616), .b(p40), .O(EX97) );
and2 gate( .a(N889), .b(EX97), .O(EX98) );
or2  gate( .a(EX92), .b(EX94), .O(EX99) );
or2  gate( .a(EX96), .b(EX99), .O(EX100) );
or2  gate( .a(EX98), .b(EX100), .O(N1055) );
nand2 gate235( .a(N625), .b(N890), .O(N1063) );
inv1 gate( .a(N622),.O(N622_NOT) );
inv1 gate( .a(N891),.O(N891_NOT));
and2 gate( .a(N622_NOT), .b(p41), .O(EX101) );
and2 gate( .a(N891_NOT), .b(EX101), .O(EX102) );
and2 gate( .a(N622), .b(p42), .O(EX103) );
and2 gate( .a(N891_NOT), .b(EX103), .O(EX104) );
and2 gate( .a(N622_NOT), .b(p43), .O(EX105) );
and2 gate( .a(N891), .b(EX105), .O(EX106) );
and2 gate( .a(N622), .b(p44), .O(EX107) );
and2 gate( .a(N891), .b(EX107), .O(EX108) );
or2  gate( .a(EX102), .b(EX104), .O(EX109) );
or2  gate( .a(EX106), .b(EX109), .O(EX110) );
or2  gate( .a(EX108), .b(EX110), .O(N1064) );
inv1 gate( .a(N655),.O(N655_NOT) );
inv1 gate( .a(N895),.O(N895_NOT));
and2 gate( .a(N655_NOT), .b(p45), .O(EX111) );
and2 gate( .a(N895_NOT), .b(EX111), .O(EX112) );
and2 gate( .a(N655), .b(p46), .O(EX113) );
and2 gate( .a(N895_NOT), .b(EX113), .O(EX114) );
and2 gate( .a(N655_NOT), .b(p47), .O(EX115) );
and2 gate( .a(N895), .b(EX115), .O(EX116) );
and2 gate( .a(N655), .b(p48), .O(EX117) );
and2 gate( .a(N895), .b(EX117), .O(EX118) );
or2  gate( .a(EX112), .b(EX114), .O(EX119) );
or2  gate( .a(EX116), .b(EX119), .O(EX120) );
or2  gate( .a(EX118), .b(EX120), .O(N1067) );
inv1 gate( .a(N652),.O(N652_NOT) );
inv1 gate( .a(N896),.O(N896_NOT));
and2 gate( .a(N652_NOT), .b(p49), .O(EX121) );
and2 gate( .a(N896_NOT), .b(EX121), .O(EX122) );
and2 gate( .a(N652), .b(p50), .O(EX123) );
and2 gate( .a(N896_NOT), .b(EX123), .O(EX124) );
and2 gate( .a(N652_NOT), .b(p51), .O(EX125) );
and2 gate( .a(N896), .b(EX125), .O(EX126) );
and2 gate( .a(N652), .b(p52), .O(EX127) );
and2 gate( .a(N896), .b(EX127), .O(EX128) );
or2  gate( .a(EX122), .b(EX124), .O(EX129) );
or2  gate( .a(EX126), .b(EX129), .O(EX130) );
or2  gate( .a(EX128), .b(EX130), .O(N1068) );
nand2 gate239( .a(N721), .b(N988), .O(N1119) );
nand2 gate240( .a(N718), .b(N989), .O(N1120) );
inv1 gate( .a(N727),.O(N727_NOT) );
inv1 gate( .a(N991),.O(N991_NOT));
and2 gate( .a(N727_NOT), .b(p53), .O(EX131) );
and2 gate( .a(N991_NOT), .b(EX131), .O(EX132) );
and2 gate( .a(N727), .b(p54), .O(EX133) );
and2 gate( .a(N991_NOT), .b(EX133), .O(EX134) );
and2 gate( .a(N727_NOT), .b(p55), .O(EX135) );
and2 gate( .a(N991), .b(EX135), .O(EX136) );
and2 gate( .a(N727), .b(p56), .O(EX137) );
and2 gate( .a(N991), .b(EX137), .O(EX138) );
or2  gate( .a(EX132), .b(EX134), .O(EX139) );
or2  gate( .a(EX136), .b(EX139), .O(EX140) );
or2  gate( .a(EX138), .b(EX140), .O(N1121) );
nand2 gate242( .a(N724), .b(N992), .O(N1122) );
inv1 gate( .a(N739),.O(N739_NOT) );
inv1 gate( .a(N1002),.O(N1002_NOT));
and2 gate( .a(N739_NOT), .b(p57), .O(EX141) );
and2 gate( .a(N1002_NOT), .b(EX141), .O(EX142) );
and2 gate( .a(N739), .b(p58), .O(EX143) );
and2 gate( .a(N1002_NOT), .b(EX143), .O(EX144) );
and2 gate( .a(N739_NOT), .b(p59), .O(EX145) );
and2 gate( .a(N1002), .b(EX145), .O(EX146) );
and2 gate( .a(N739), .b(p60), .O(EX147) );
and2 gate( .a(N1002), .b(EX147), .O(EX148) );
or2  gate( .a(EX142), .b(EX144), .O(EX149) );
or2  gate( .a(EX146), .b(EX149), .O(EX150) );
or2  gate( .a(EX148), .b(EX150), .O(N1128) );
nand2 gate244( .a(N736), .b(N1003), .O(N1129) );
nand2 gate245( .a(N745), .b(N1005), .O(N1130) );
nand2 gate246( .a(N742), .b(N1006), .O(N1131) );
nand2 gate247( .a(N751), .b(N1008), .O(N1132) );
inv1 gate( .a(N748),.O(N748_NOT) );
inv1 gate( .a(N1009),.O(N1009_NOT));
and2 gate( .a(N748_NOT), .b(p61), .O(EX151) );
and2 gate( .a(N1009_NOT), .b(EX151), .O(EX152) );
and2 gate( .a(N748), .b(p62), .O(EX153) );
and2 gate( .a(N1009_NOT), .b(EX153), .O(EX154) );
and2 gate( .a(N748_NOT), .b(p63), .O(EX155) );
and2 gate( .a(N1009), .b(EX155), .O(EX156) );
and2 gate( .a(N748), .b(p64), .O(EX157) );
and2 gate( .a(N1009), .b(EX157), .O(EX158) );
or2  gate( .a(EX152), .b(EX154), .O(EX159) );
or2  gate( .a(EX156), .b(EX159), .O(EX160) );
or2  gate( .a(EX158), .b(EX160), .O(N1133) );
inv1 gate249( .a(N939), .O(N1148) );
inv1 gate250( .a(N935), .O(N1149) );
inv1 gate( .a(N1054),.O(N1054_NOT) );
inv1 gate( .a(N1055),.O(N1055_NOT));
and2 gate( .a(N1054_NOT), .b(p65), .O(EX161) );
and2 gate( .a(N1055_NOT), .b(EX161), .O(EX162) );
and2 gate( .a(N1054), .b(p66), .O(EX163) );
and2 gate( .a(N1055_NOT), .b(EX163), .O(EX164) );
and2 gate( .a(N1054_NOT), .b(p67), .O(EX165) );
and2 gate( .a(N1055), .b(EX165), .O(EX166) );
and2 gate( .a(N1054), .b(p68), .O(EX167) );
and2 gate( .a(N1055), .b(EX167), .O(EX168) );
or2  gate( .a(EX162), .b(EX164), .O(EX169) );
or2  gate( .a(EX166), .b(EX169), .O(EX170) );
or2  gate( .a(EX168), .b(EX170), .O(N1150) );
inv1 gate252( .a(N943), .O(N1151) );
inv1 gate253( .a(N947), .O(N1152) );
inv1 gate254( .a(N955), .O(N1153) );
inv1 gate255( .a(N951), .O(N1154) );
inv1 gate256( .a(N962), .O(N1155) );
inv1 gate257( .a(N969), .O(N1156) );
inv1 gate258( .a(N977), .O(N1157) );
nand2 gate259( .a(N1063), .b(N1064), .O(N1158) );
inv1 gate260( .a(N985), .O(N1159) );
inv1 gate( .a(N985),.O(N985_NOT) );
inv1 gate( .a(N892),.O(N892_NOT));
and2 gate( .a(N985_NOT), .b(p69), .O(EX171) );
and2 gate( .a(N892_NOT), .b(EX171), .O(EX172) );
and2 gate( .a(N985), .b(p70), .O(EX173) );
and2 gate( .a(N892_NOT), .b(EX173), .O(EX174) );
and2 gate( .a(N985_NOT), .b(p71), .O(EX175) );
and2 gate( .a(N892), .b(EX175), .O(EX176) );
and2 gate( .a(N985), .b(p72), .O(EX177) );
and2 gate( .a(N892), .b(EX177), .O(EX178) );
or2  gate( .a(EX172), .b(EX174), .O(EX179) );
or2  gate( .a(EX176), .b(EX179), .O(EX180) );
or2  gate( .a(EX178), .b(EX180), .O(N1160) );
inv1 gate262( .a(N998), .O(N1161) );
nand2 gate263( .a(N1067), .b(N1068), .O(N1162) );
inv1 gate264( .a(N899), .O(N1163) );
buf1 gate265( .a(N899), .O(N1164) );
inv1 gate266( .a(N903), .O(N1167) );
buf1 gate267( .a(N903), .O(N1168) );
nand2 gate268( .a(N921), .b(N923), .O(N1171) );
inv1 gate( .a(N922),.O(N922_NOT) );
inv1 gate( .a(N923),.O(N923_NOT));
and2 gate( .a(N922_NOT), .b(p73), .O(EX181) );
and2 gate( .a(N923_NOT), .b(EX181), .O(EX182) );
and2 gate( .a(N922), .b(p74), .O(EX183) );
and2 gate( .a(N923_NOT), .b(EX183), .O(EX184) );
and2 gate( .a(N922_NOT), .b(p75), .O(EX185) );
and2 gate( .a(N923), .b(EX185), .O(EX186) );
and2 gate( .a(N922), .b(p76), .O(EX187) );
and2 gate( .a(N923), .b(EX187), .O(EX188) );
or2  gate( .a(EX182), .b(EX184), .O(EX189) );
or2  gate( .a(EX186), .b(EX189), .O(EX190) );
or2  gate( .a(EX188), .b(EX190), .O(N1188) );
inv1 gate270( .a(N1010), .O(N1205) );
nand2 gate271( .a(N1010), .b(N938), .O(N1206) );
inv1 gate272( .a(N1013), .O(N1207) );
nand2 gate273( .a(N1013), .b(N942), .O(N1208) );
inv1 gate274( .a(N1016), .O(N1209) );
nand2 gate275( .a(N1016), .b(N946), .O(N1210) );
inv1 gate276( .a(N1019), .O(N1211) );
nand2 gate277( .a(N1019), .b(N950), .O(N1212) );
inv1 gate278( .a(N1022), .O(N1213) );
nand2 gate279( .a(N1022), .b(N954), .O(N1214) );
inv1 gate280( .a(N1025), .O(N1215) );
nand2 gate281( .a(N1025), .b(N958), .O(N1216) );
inv1 gate282( .a(N1028), .O(N1217) );
inv1 gate283( .a(N959), .O(N1218) );
inv1 gate284( .a(N1031), .O(N1219) );
inv1 gate285( .a(N1034), .O(N1220) );
nand2 gate286( .a(N1034), .b(N968), .O(N1221) );
inv1 gate287( .a(N965), .O(N1222) );
inv1 gate288( .a(N1037), .O(N1223) );
nand2 gate289( .a(N1037), .b(N972), .O(N1224) );
inv1 gate290( .a(N1040), .O(N1225) );
nand2 gate291( .a(N1040), .b(N976), .O(N1226) );
inv1 gate292( .a(N973), .O(N1227) );
inv1 gate293( .a(N1043), .O(N1228) );
nand2 gate294( .a(N1043), .b(N980), .O(N1229) );
inv1 gate295( .a(N981), .O(N1230) );
inv1 gate( .a(N981),.O(N981_NOT) );
inv1 gate( .a(N984),.O(N984_NOT));
and2 gate( .a(N981_NOT), .b(p77), .O(EX191) );
and2 gate( .a(N984_NOT), .b(EX191), .O(EX192) );
and2 gate( .a(N981), .b(p78), .O(EX193) );
and2 gate( .a(N984_NOT), .b(EX193), .O(EX194) );
and2 gate( .a(N981_NOT), .b(p79), .O(EX195) );
and2 gate( .a(N984), .b(EX195), .O(EX196) );
and2 gate( .a(N981), .b(p80), .O(EX197) );
and2 gate( .a(N984), .b(EX197), .O(EX198) );
or2  gate( .a(EX192), .b(EX194), .O(EX199) );
or2  gate( .a(EX196), .b(EX199), .O(EX200) );
or2  gate( .a(EX198), .b(EX200), .O(N1231) );
nand2 gate297( .a(N1119), .b(N1120), .O(N1232) );
nand2 gate298( .a(N1121), .b(N1122), .O(N1235) );
inv1 gate299( .a(N1046), .O(N1238) );
nand2 gate300( .a(N1046), .b(N997), .O(N1239) );
inv1 gate301( .a(N994), .O(N1240) );
inv1 gate302( .a(N1049), .O(N1241) );
inv1 gate( .a(N1049),.O(N1049_NOT) );
inv1 gate( .a(N1001),.O(N1001_NOT));
and2 gate( .a(N1049_NOT), .b(p81), .O(EX201) );
and2 gate( .a(N1001_NOT), .b(EX201), .O(EX202) );
and2 gate( .a(N1049), .b(p82), .O(EX203) );
and2 gate( .a(N1001_NOT), .b(EX203), .O(EX204) );
and2 gate( .a(N1049_NOT), .b(p83), .O(EX205) );
and2 gate( .a(N1001), .b(EX205), .O(EX206) );
and2 gate( .a(N1049), .b(p84), .O(EX207) );
and2 gate( .a(N1001), .b(EX207), .O(EX208) );
or2  gate( .a(EX202), .b(EX204), .O(EX209) );
or2  gate( .a(EX206), .b(EX209), .O(EX210) );
or2  gate( .a(EX208), .b(EX210), .O(N1242) );
nand2 gate304( .a(N1128), .b(N1129), .O(N1243) );
nand2 gate305( .a(N1130), .b(N1131), .O(N1246) );
inv1 gate( .a(N1132),.O(N1132_NOT) );
inv1 gate( .a(N1133),.O(N1133_NOT));
and2 gate( .a(N1132_NOT), .b(p85), .O(EX211) );
and2 gate( .a(N1133_NOT), .b(EX211), .O(EX212) );
and2 gate( .a(N1132), .b(p86), .O(EX213) );
and2 gate( .a(N1133_NOT), .b(EX213), .O(EX214) );
and2 gate( .a(N1132_NOT), .b(p87), .O(EX215) );
and2 gate( .a(N1133), .b(EX215), .O(EX216) );
and2 gate( .a(N1132), .b(p88), .O(EX217) );
and2 gate( .a(N1133), .b(EX217), .O(EX218) );
or2  gate( .a(EX212), .b(EX214), .O(EX219) );
or2  gate( .a(EX216), .b(EX219), .O(EX220) );
or2  gate( .a(EX218), .b(EX220), .O(N1249) );
buf1 gate307( .a(N907), .O(N1252) );
buf1 gate308( .a(N907), .O(N1255) );
buf1 gate309( .a(N910), .O(N1258) );
buf1 gate310( .a(N910), .O(N1261) );
inv1 gate311( .a(N1150), .O(N1264) );
nand2 gate312( .a(N631), .b(N1159), .O(N1267) );
nand2 gate313( .a(N688), .b(N1205), .O(N1309) );
nand2 gate314( .a(N691), .b(N1207), .O(N1310) );
nand2 gate315( .a(N694), .b(N1209), .O(N1311) );
nand2 gate316( .a(N697), .b(N1211), .O(N1312) );
nand2 gate317( .a(N700), .b(N1213), .O(N1313) );
nand2 gate318( .a(N703), .b(N1215), .O(N1314) );
nand2 gate319( .a(N706), .b(N1220), .O(N1315) );
inv1 gate( .a(N709),.O(N709_NOT) );
inv1 gate( .a(N1223),.O(N1223_NOT));
and2 gate( .a(N709_NOT), .b(p89), .O(EX221) );
and2 gate( .a(N1223_NOT), .b(EX221), .O(EX222) );
and2 gate( .a(N709), .b(p90), .O(EX223) );
and2 gate( .a(N1223_NOT), .b(EX223), .O(EX224) );
and2 gate( .a(N709_NOT), .b(p91), .O(EX225) );
and2 gate( .a(N1223), .b(EX225), .O(EX226) );
and2 gate( .a(N709), .b(p92), .O(EX227) );
and2 gate( .a(N1223), .b(EX227), .O(EX228) );
or2  gate( .a(EX222), .b(EX224), .O(EX229) );
or2  gate( .a(EX226), .b(EX229), .O(EX230) );
or2  gate( .a(EX228), .b(EX230), .O(N1316) );
inv1 gate( .a(N712),.O(N712_NOT) );
inv1 gate( .a(N1225),.O(N1225_NOT));
and2 gate( .a(N712_NOT), .b(p93), .O(EX231) );
and2 gate( .a(N1225_NOT), .b(EX231), .O(EX232) );
and2 gate( .a(N712), .b(p94), .O(EX233) );
and2 gate( .a(N1225_NOT), .b(EX233), .O(EX234) );
and2 gate( .a(N712_NOT), .b(p95), .O(EX235) );
and2 gate( .a(N1225), .b(EX235), .O(EX236) );
and2 gate( .a(N712), .b(p96), .O(EX237) );
and2 gate( .a(N1225), .b(EX237), .O(EX238) );
or2  gate( .a(EX232), .b(EX234), .O(EX239) );
or2  gate( .a(EX236), .b(EX239), .O(EX240) );
or2  gate( .a(EX238), .b(EX240), .O(N1317) );
nand2 gate322( .a(N715), .b(N1228), .O(N1318) );
inv1 gate323( .a(N1158), .O(N1319) );
inv1 gate( .a(N628),.O(N628_NOT) );
inv1 gate( .a(N1230),.O(N1230_NOT));
and2 gate( .a(N628_NOT), .b(p97), .O(EX241) );
and2 gate( .a(N1230_NOT), .b(EX241), .O(EX242) );
and2 gate( .a(N628), .b(p98), .O(EX243) );
and2 gate( .a(N1230_NOT), .b(EX243), .O(EX244) );
and2 gate( .a(N628_NOT), .b(p99), .O(EX245) );
and2 gate( .a(N1230), .b(EX245), .O(EX246) );
and2 gate( .a(N628), .b(p100), .O(EX247) );
and2 gate( .a(N1230), .b(EX247), .O(EX248) );
or2  gate( .a(EX242), .b(EX244), .O(EX249) );
or2  gate( .a(EX246), .b(EX249), .O(EX250) );
or2  gate( .a(EX248), .b(EX250), .O(N1322) );
inv1 gate( .a(N730),.O(N730_NOT) );
inv1 gate( .a(N1238),.O(N1238_NOT));
and2 gate( .a(N730_NOT), .b(p101), .O(EX251) );
and2 gate( .a(N1238_NOT), .b(EX251), .O(EX252) );
and2 gate( .a(N730), .b(p102), .O(EX253) );
and2 gate( .a(N1238_NOT), .b(EX253), .O(EX254) );
and2 gate( .a(N730_NOT), .b(p103), .O(EX255) );
and2 gate( .a(N1238), .b(EX255), .O(EX256) );
and2 gate( .a(N730), .b(p104), .O(EX257) );
and2 gate( .a(N1238), .b(EX257), .O(EX258) );
or2  gate( .a(EX252), .b(EX254), .O(EX259) );
or2  gate( .a(EX256), .b(EX259), .O(EX260) );
or2  gate( .a(EX258), .b(EX260), .O(N1327) );
nand2 gate326( .a(N733), .b(N1241), .O(N1328) );
inv1 gate327( .a(N1162), .O(N1334) );
inv1 gate( .a(N1267),.O(N1267_NOT) );
inv1 gate( .a(N1160),.O(N1160_NOT));
and2 gate( .a(N1267_NOT), .b(p105), .O(EX261) );
and2 gate( .a(N1160_NOT), .b(EX261), .O(EX262) );
and2 gate( .a(N1267), .b(p106), .O(EX263) );
and2 gate( .a(N1160_NOT), .b(EX263), .O(EX264) );
and2 gate( .a(N1267_NOT), .b(p107), .O(EX265) );
and2 gate( .a(N1160), .b(EX265), .O(EX266) );
and2 gate( .a(N1267), .b(p108), .O(EX267) );
and2 gate( .a(N1160), .b(EX267), .O(EX268) );
or2  gate( .a(EX262), .b(EX264), .O(EX269) );
or2  gate( .a(EX266), .b(EX269), .O(EX270) );
or2  gate( .a(EX268), .b(EX270), .O(N1344) );
nand2 gate329( .a(N1249), .b(N894), .O(N1345) );
inv1 gate330( .a(N1249), .O(N1346) );
inv1 gate331( .a(N1255), .O(N1348) );
inv1 gate332( .a(N1252), .O(N1349) );
inv1 gate333( .a(N1261), .O(N1350) );
inv1 gate334( .a(N1258), .O(N1351) );
nand2 gate335( .a(N1309), .b(N1206), .O(N1352) );
nand2 gate336( .a(N1310), .b(N1208), .O(N1355) );
inv1 gate( .a(N1311),.O(N1311_NOT) );
inv1 gate( .a(N1210),.O(N1210_NOT));
and2 gate( .a(N1311_NOT), .b(p109), .O(EX271) );
and2 gate( .a(N1210_NOT), .b(EX271), .O(EX272) );
and2 gate( .a(N1311), .b(p110), .O(EX273) );
and2 gate( .a(N1210_NOT), .b(EX273), .O(EX274) );
and2 gate( .a(N1311_NOT), .b(p111), .O(EX275) );
and2 gate( .a(N1210), .b(EX275), .O(EX276) );
and2 gate( .a(N1311), .b(p112), .O(EX277) );
and2 gate( .a(N1210), .b(EX277), .O(EX278) );
or2  gate( .a(EX272), .b(EX274), .O(EX279) );
or2  gate( .a(EX276), .b(EX279), .O(EX280) );
or2  gate( .a(EX278), .b(EX280), .O(N1358) );
inv1 gate( .a(N1312),.O(N1312_NOT) );
inv1 gate( .a(N1212),.O(N1212_NOT));
and2 gate( .a(N1312_NOT), .b(p113), .O(EX281) );
and2 gate( .a(N1212_NOT), .b(EX281), .O(EX282) );
and2 gate( .a(N1312), .b(p114), .O(EX283) );
and2 gate( .a(N1212_NOT), .b(EX283), .O(EX284) );
and2 gate( .a(N1312_NOT), .b(p115), .O(EX285) );
and2 gate( .a(N1212), .b(EX285), .O(EX286) );
and2 gate( .a(N1312), .b(p116), .O(EX287) );
and2 gate( .a(N1212), .b(EX287), .O(EX288) );
or2  gate( .a(EX282), .b(EX284), .O(EX289) );
or2  gate( .a(EX286), .b(EX289), .O(EX290) );
or2  gate( .a(EX288), .b(EX290), .O(N1361) );
nand2 gate339( .a(N1313), .b(N1214), .O(N1364) );
nand2 gate340( .a(N1314), .b(N1216), .O(N1367) );
nand2 gate341( .a(N1315), .b(N1221), .O(N1370) );
nand2 gate342( .a(N1316), .b(N1224), .O(N1373) );
inv1 gate( .a(N1317),.O(N1317_NOT) );
inv1 gate( .a(N1226),.O(N1226_NOT));
and2 gate( .a(N1317_NOT), .b(p117), .O(EX291) );
and2 gate( .a(N1226_NOT), .b(EX291), .O(EX292) );
and2 gate( .a(N1317), .b(p118), .O(EX293) );
and2 gate( .a(N1226_NOT), .b(EX293), .O(EX294) );
and2 gate( .a(N1317_NOT), .b(p119), .O(EX295) );
and2 gate( .a(N1226), .b(EX295), .O(EX296) );
and2 gate( .a(N1317), .b(p120), .O(EX297) );
and2 gate( .a(N1226), .b(EX297), .O(EX298) );
or2  gate( .a(EX292), .b(EX294), .O(EX299) );
or2  gate( .a(EX296), .b(EX299), .O(EX300) );
or2  gate( .a(EX298), .b(EX300), .O(N1376) );
nand2 gate344( .a(N1318), .b(N1229), .O(N1379) );
inv1 gate( .a(N1322),.O(N1322_NOT) );
inv1 gate( .a(N1231),.O(N1231_NOT));
and2 gate( .a(N1322_NOT), .b(p121), .O(EX301) );
and2 gate( .a(N1231_NOT), .b(EX301), .O(EX302) );
and2 gate( .a(N1322), .b(p122), .O(EX303) );
and2 gate( .a(N1231_NOT), .b(EX303), .O(EX304) );
and2 gate( .a(N1322_NOT), .b(p123), .O(EX305) );
and2 gate( .a(N1231), .b(EX305), .O(EX306) );
and2 gate( .a(N1322), .b(p124), .O(EX307) );
and2 gate( .a(N1231), .b(EX307), .O(EX308) );
or2  gate( .a(EX302), .b(EX304), .O(EX309) );
or2  gate( .a(EX306), .b(EX309), .O(EX310) );
or2  gate( .a(EX308), .b(EX310), .O(N1383) );
inv1 gate346( .a(N1232), .O(N1386) );
inv1 gate( .a(N1232),.O(N1232_NOT) );
inv1 gate( .a(N990),.O(N990_NOT));
and2 gate( .a(N1232_NOT), .b(p125), .O(EX311) );
and2 gate( .a(N990_NOT), .b(EX311), .O(EX312) );
and2 gate( .a(N1232), .b(p126), .O(EX313) );
and2 gate( .a(N990_NOT), .b(EX313), .O(EX314) );
and2 gate( .a(N1232_NOT), .b(p127), .O(EX315) );
and2 gate( .a(N990), .b(EX315), .O(EX316) );
and2 gate( .a(N1232), .b(p128), .O(EX317) );
and2 gate( .a(N990), .b(EX317), .O(EX318) );
or2  gate( .a(EX312), .b(EX314), .O(EX319) );
or2  gate( .a(EX316), .b(EX319), .O(EX320) );
or2  gate( .a(EX318), .b(EX320), .O(N1387) );
inv1 gate348( .a(N1235), .O(N1388) );
inv1 gate( .a(N1235),.O(N1235_NOT) );
inv1 gate( .a(N993),.O(N993_NOT));
and2 gate( .a(N1235_NOT), .b(p129), .O(EX321) );
and2 gate( .a(N993_NOT), .b(EX321), .O(EX322) );
and2 gate( .a(N1235), .b(p130), .O(EX323) );
and2 gate( .a(N993_NOT), .b(EX323), .O(EX324) );
and2 gate( .a(N1235_NOT), .b(p131), .O(EX325) );
and2 gate( .a(N993), .b(EX325), .O(EX326) );
and2 gate( .a(N1235), .b(p132), .O(EX327) );
and2 gate( .a(N993), .b(EX327), .O(EX328) );
or2  gate( .a(EX322), .b(EX324), .O(EX329) );
or2  gate( .a(EX326), .b(EX329), .O(EX330) );
or2  gate( .a(EX328), .b(EX330), .O(N1389) );
nand2 gate350( .a(N1327), .b(N1239), .O(N1390) );
nand2 gate351( .a(N1328), .b(N1242), .O(N1393) );
inv1 gate352( .a(N1243), .O(N1396) );
nand2 gate353( .a(N1243), .b(N1004), .O(N1397) );
inv1 gate354( .a(N1246), .O(N1398) );
nand2 gate355( .a(N1246), .b(N1007), .O(N1399) );
inv1 gate356( .a(N1319), .O(N1409) );
inv1 gate( .a(N649),.O(N649_NOT) );
inv1 gate( .a(N1346),.O(N1346_NOT));
and2 gate( .a(N649_NOT), .b(p133), .O(EX331) );
and2 gate( .a(N1346_NOT), .b(EX331), .O(EX332) );
and2 gate( .a(N649), .b(p134), .O(EX333) );
and2 gate( .a(N1346_NOT), .b(EX333), .O(EX334) );
and2 gate( .a(N649_NOT), .b(p135), .O(EX335) );
and2 gate( .a(N1346), .b(EX335), .O(EX336) );
and2 gate( .a(N649), .b(p136), .O(EX337) );
and2 gate( .a(N1346), .b(EX337), .O(EX338) );
or2  gate( .a(EX332), .b(EX334), .O(EX339) );
or2  gate( .a(EX336), .b(EX339), .O(EX340) );
or2  gate( .a(EX338), .b(EX340), .O(N1412) );
inv1 gate358( .a(N1334), .O(N1413) );
buf1 gate359( .a(N1264), .O(N1416) );
buf1 gate360( .a(N1264), .O(N1419) );
nand2 gate361( .a(N634), .b(N1386), .O(N1433) );
inv1 gate( .a(N637),.O(N637_NOT) );
inv1 gate( .a(N1388),.O(N1388_NOT));
and2 gate( .a(N637_NOT), .b(p137), .O(EX341) );
and2 gate( .a(N1388_NOT), .b(EX341), .O(EX342) );
and2 gate( .a(N637), .b(p138), .O(EX343) );
and2 gate( .a(N1388_NOT), .b(EX343), .O(EX344) );
and2 gate( .a(N637_NOT), .b(p139), .O(EX345) );
and2 gate( .a(N1388), .b(EX345), .O(EX346) );
and2 gate( .a(N637), .b(p140), .O(EX347) );
and2 gate( .a(N1388), .b(EX347), .O(EX348) );
or2  gate( .a(EX342), .b(EX344), .O(EX349) );
or2  gate( .a(EX346), .b(EX349), .O(EX350) );
or2  gate( .a(EX348), .b(EX350), .O(N1434) );
nand2 gate363( .a(N640), .b(N1396), .O(N1438) );
nand2 gate364( .a(N646), .b(N1398), .O(N1439) );
inv1 gate365( .a(N1344), .O(N1440) );
nand2 gate366( .a(N1355), .b(N1148), .O(N1443) );
inv1 gate367( .a(N1355), .O(N1444) );
inv1 gate( .a(N1352),.O(N1352_NOT) );
inv1 gate( .a(N1149),.O(N1149_NOT));
and2 gate( .a(N1352_NOT), .b(p141), .O(EX351) );
and2 gate( .a(N1149_NOT), .b(EX351), .O(EX352) );
and2 gate( .a(N1352), .b(p142), .O(EX353) );
and2 gate( .a(N1149_NOT), .b(EX353), .O(EX354) );
and2 gate( .a(N1352_NOT), .b(p143), .O(EX355) );
and2 gate( .a(N1149), .b(EX355), .O(EX356) );
and2 gate( .a(N1352), .b(p144), .O(EX357) );
and2 gate( .a(N1149), .b(EX357), .O(EX358) );
or2  gate( .a(EX352), .b(EX354), .O(EX359) );
or2  gate( .a(EX356), .b(EX359), .O(EX360) );
or2  gate( .a(EX358), .b(EX360), .O(N1445) );
inv1 gate369( .a(N1352), .O(N1446) );
nand2 gate370( .a(N1358), .b(N1151), .O(N1447) );
inv1 gate371( .a(N1358), .O(N1448) );
inv1 gate( .a(N1361),.O(N1361_NOT) );
inv1 gate( .a(N1152),.O(N1152_NOT));
and2 gate( .a(N1361_NOT), .b(p145), .O(EX361) );
and2 gate( .a(N1152_NOT), .b(EX361), .O(EX362) );
and2 gate( .a(N1361), .b(p146), .O(EX363) );
and2 gate( .a(N1152_NOT), .b(EX363), .O(EX364) );
and2 gate( .a(N1361_NOT), .b(p147), .O(EX365) );
and2 gate( .a(N1152), .b(EX365), .O(EX366) );
and2 gate( .a(N1361), .b(p148), .O(EX367) );
and2 gate( .a(N1152), .b(EX367), .O(EX368) );
or2  gate( .a(EX362), .b(EX364), .O(EX369) );
or2  gate( .a(EX366), .b(EX369), .O(EX370) );
or2  gate( .a(EX368), .b(EX370), .O(N1451) );
inv1 gate373( .a(N1361), .O(N1452) );
nand2 gate374( .a(N1367), .b(N1153), .O(N1453) );
inv1 gate375( .a(N1367), .O(N1454) );
nand2 gate376( .a(N1364), .b(N1154), .O(N1455) );
inv1 gate377( .a(N1364), .O(N1456) );
nand2 gate378( .a(N1373), .b(N1156), .O(N1457) );
inv1 gate379( .a(N1373), .O(N1458) );
inv1 gate( .a(N1379),.O(N1379_NOT) );
inv1 gate( .a(N1157),.O(N1157_NOT));
and2 gate( .a(N1379_NOT), .b(p149), .O(EX371) );
and2 gate( .a(N1157_NOT), .b(EX371), .O(EX372) );
and2 gate( .a(N1379), .b(p150), .O(EX373) );
and2 gate( .a(N1157_NOT), .b(EX373), .O(EX374) );
and2 gate( .a(N1379_NOT), .b(p151), .O(EX375) );
and2 gate( .a(N1157), .b(EX375), .O(EX376) );
and2 gate( .a(N1379), .b(p152), .O(EX377) );
and2 gate( .a(N1157), .b(EX377), .O(EX378) );
or2  gate( .a(EX372), .b(EX374), .O(EX379) );
or2  gate( .a(EX376), .b(EX379), .O(EX380) );
or2  gate( .a(EX378), .b(EX380), .O(N1459) );
inv1 gate381( .a(N1379), .O(N1460) );
inv1 gate382( .a(N1383), .O(N1461) );
nand2 gate383( .a(N1393), .b(N1161), .O(N1462) );
inv1 gate384( .a(N1393), .O(N1463) );
nand2 gate385( .a(N1345), .b(N1412), .O(N1464) );
inv1 gate386( .a(N1370), .O(N1468) );
nand2 gate387( .a(N1370), .b(N1222), .O(N1469) );
inv1 gate388( .a(N1376), .O(N1470) );
inv1 gate( .a(N1376),.O(N1376_NOT) );
inv1 gate( .a(N1227),.O(N1227_NOT));
and2 gate( .a(N1376_NOT), .b(p153), .O(EX381) );
and2 gate( .a(N1227_NOT), .b(EX381), .O(EX382) );
and2 gate( .a(N1376), .b(p154), .O(EX383) );
and2 gate( .a(N1227_NOT), .b(EX383), .O(EX384) );
and2 gate( .a(N1376_NOT), .b(p155), .O(EX385) );
and2 gate( .a(N1227), .b(EX385), .O(EX386) );
and2 gate( .a(N1376), .b(p156), .O(EX387) );
and2 gate( .a(N1227), .b(EX387), .O(EX388) );
or2  gate( .a(EX382), .b(EX384), .O(EX389) );
or2  gate( .a(EX386), .b(EX389), .O(EX390) );
or2  gate( .a(EX388), .b(EX390), .O(N1471) );
nand2 gate390( .a(N1387), .b(N1433), .O(N1472) );
inv1 gate391( .a(N1390), .O(N1475) );
nand2 gate392( .a(N1390), .b(N1240), .O(N1476) );
nand2 gate393( .a(N1389), .b(N1434), .O(N1478) );
nand2 gate394( .a(N1399), .b(N1439), .O(N1481) );
inv1 gate( .a(N1397),.O(N1397_NOT) );
inv1 gate( .a(N1438),.O(N1438_NOT));
and2 gate( .a(N1397_NOT), .b(p157), .O(EX391) );
and2 gate( .a(N1438_NOT), .b(EX391), .O(EX392) );
and2 gate( .a(N1397), .b(p158), .O(EX393) );
and2 gate( .a(N1438_NOT), .b(EX393), .O(EX394) );
and2 gate( .a(N1397_NOT), .b(p159), .O(EX395) );
and2 gate( .a(N1438), .b(EX395), .O(EX396) );
and2 gate( .a(N1397), .b(p160), .O(EX397) );
and2 gate( .a(N1438), .b(EX397), .O(EX398) );
or2  gate( .a(EX392), .b(EX394), .O(EX399) );
or2  gate( .a(EX396), .b(EX399), .O(EX400) );
or2  gate( .a(EX398), .b(EX400), .O(N1484) );
inv1 gate( .a(N939),.O(N939_NOT) );
inv1 gate( .a(N1444),.O(N1444_NOT));
and2 gate( .a(N939_NOT), .b(p161), .O(EX401) );
and2 gate( .a(N1444_NOT), .b(EX401), .O(EX402) );
and2 gate( .a(N939), .b(p162), .O(EX403) );
and2 gate( .a(N1444_NOT), .b(EX403), .O(EX404) );
and2 gate( .a(N939_NOT), .b(p163), .O(EX405) );
and2 gate( .a(N1444), .b(EX405), .O(EX406) );
and2 gate( .a(N939), .b(p164), .O(EX407) );
and2 gate( .a(N1444), .b(EX407), .O(EX408) );
or2  gate( .a(EX402), .b(EX404), .O(EX409) );
or2  gate( .a(EX406), .b(EX409), .O(EX410) );
or2  gate( .a(EX408), .b(EX410), .O(N1487) );
inv1 gate( .a(N935),.O(N935_NOT) );
inv1 gate( .a(N1446),.O(N1446_NOT));
and2 gate( .a(N935_NOT), .b(p165), .O(EX411) );
and2 gate( .a(N1446_NOT), .b(EX411), .O(EX412) );
and2 gate( .a(N935), .b(p166), .O(EX413) );
and2 gate( .a(N1446_NOT), .b(EX413), .O(EX414) );
and2 gate( .a(N935_NOT), .b(p167), .O(EX415) );
and2 gate( .a(N1446), .b(EX415), .O(EX416) );
and2 gate( .a(N935), .b(p168), .O(EX417) );
and2 gate( .a(N1446), .b(EX417), .O(EX418) );
or2  gate( .a(EX412), .b(EX414), .O(EX419) );
or2  gate( .a(EX416), .b(EX419), .O(EX420) );
or2  gate( .a(EX418), .b(EX420), .O(N1488) );
nand2 gate398( .a(N943), .b(N1448), .O(N1489) );
inv1 gate399( .a(N1419), .O(N1490) );
inv1 gate400( .a(N1416), .O(N1491) );
nand2 gate401( .a(N947), .b(N1452), .O(N1492) );
nand2 gate402( .a(N955), .b(N1454), .O(N1493) );
nand2 gate403( .a(N951), .b(N1456), .O(N1494) );
nand2 gate404( .a(N969), .b(N1458), .O(N1495) );
nand2 gate405( .a(N977), .b(N1460), .O(N1496) );
inv1 gate( .a(N998),.O(N998_NOT) );
inv1 gate( .a(N1463),.O(N1463_NOT));
and2 gate( .a(N998_NOT), .b(p169), .O(EX421) );
and2 gate( .a(N1463_NOT), .b(EX421), .O(EX422) );
and2 gate( .a(N998), .b(p170), .O(EX423) );
and2 gate( .a(N1463_NOT), .b(EX423), .O(EX424) );
and2 gate( .a(N998_NOT), .b(p171), .O(EX425) );
and2 gate( .a(N1463), .b(EX425), .O(EX426) );
and2 gate( .a(N998), .b(p172), .O(EX427) );
and2 gate( .a(N1463), .b(EX427), .O(EX428) );
or2  gate( .a(EX422), .b(EX424), .O(EX429) );
or2  gate( .a(EX426), .b(EX429), .O(EX430) );
or2  gate( .a(EX428), .b(EX430), .O(N1498) );
inv1 gate407( .a(N1440), .O(N1499) );
inv1 gate( .a(N965),.O(N965_NOT) );
inv1 gate( .a(N1468),.O(N1468_NOT));
and2 gate( .a(N965_NOT), .b(p173), .O(EX431) );
and2 gate( .a(N1468_NOT), .b(EX431), .O(EX432) );
and2 gate( .a(N965), .b(p174), .O(EX433) );
and2 gate( .a(N1468_NOT), .b(EX433), .O(EX434) );
and2 gate( .a(N965_NOT), .b(p175), .O(EX435) );
and2 gate( .a(N1468), .b(EX435), .O(EX436) );
and2 gate( .a(N965), .b(p176), .O(EX437) );
and2 gate( .a(N1468), .b(EX437), .O(EX438) );
or2  gate( .a(EX432), .b(EX434), .O(EX439) );
or2  gate( .a(EX436), .b(EX439), .O(EX440) );
or2  gate( .a(EX438), .b(EX440), .O(N1500) );
nand2 gate409( .a(N973), .b(N1470), .O(N1501) );
nand2 gate410( .a(N994), .b(N1475), .O(N1504) );
inv1 gate411( .a(N1464), .O(N1510) );
nand2 gate412( .a(N1443), .b(N1487), .O(N1513) );
nand2 gate413( .a(N1445), .b(N1488), .O(N1514) );
nand2 gate414( .a(N1447), .b(N1489), .O(N1517) );
nand2 gate415( .a(N1451), .b(N1492), .O(N1520) );
inv1 gate( .a(N1453),.O(N1453_NOT) );
inv1 gate( .a(N1493),.O(N1493_NOT));
and2 gate( .a(N1453_NOT), .b(p177), .O(EX441) );
and2 gate( .a(N1493_NOT), .b(EX441), .O(EX442) );
and2 gate( .a(N1453), .b(p178), .O(EX443) );
and2 gate( .a(N1493_NOT), .b(EX443), .O(EX444) );
and2 gate( .a(N1453_NOT), .b(p179), .O(EX445) );
and2 gate( .a(N1493), .b(EX445), .O(EX446) );
and2 gate( .a(N1453), .b(p180), .O(EX447) );
and2 gate( .a(N1493), .b(EX447), .O(EX448) );
or2  gate( .a(EX442), .b(EX444), .O(EX449) );
or2  gate( .a(EX446), .b(EX449), .O(EX450) );
or2  gate( .a(EX448), .b(EX450), .O(N1521) );
inv1 gate( .a(N1455),.O(N1455_NOT) );
inv1 gate( .a(N1494),.O(N1494_NOT));
and2 gate( .a(N1455_NOT), .b(p181), .O(EX451) );
and2 gate( .a(N1494_NOT), .b(EX451), .O(EX452) );
and2 gate( .a(N1455), .b(p182), .O(EX453) );
and2 gate( .a(N1494_NOT), .b(EX453), .O(EX454) );
and2 gate( .a(N1455_NOT), .b(p183), .O(EX455) );
and2 gate( .a(N1494), .b(EX455), .O(EX456) );
and2 gate( .a(N1455), .b(p184), .O(EX457) );
and2 gate( .a(N1494), .b(EX457), .O(EX458) );
or2  gate( .a(EX452), .b(EX454), .O(EX459) );
or2  gate( .a(EX456), .b(EX459), .O(EX460) );
or2  gate( .a(EX458), .b(EX460), .O(N1522) );
nand2 gate418( .a(N1457), .b(N1495), .O(N1526) );
nand2 gate419( .a(N1459), .b(N1496), .O(N1527) );
inv1 gate420( .a(N1472), .O(N1528) );
nand2 gate421( .a(N1462), .b(N1498), .O(N1529) );
inv1 gate422( .a(N1478), .O(N1530) );
inv1 gate423( .a(N1481), .O(N1531) );
inv1 gate424( .a(N1484), .O(N1532) );
nand2 gate425( .a(N1471), .b(N1501), .O(N1534) );
nand2 gate426( .a(N1469), .b(N1500), .O(N1537) );
inv1 gate( .a(N1476),.O(N1476_NOT) );
inv1 gate( .a(N1504),.O(N1504_NOT));
and2 gate( .a(N1476_NOT), .b(p185), .O(EX461) );
and2 gate( .a(N1504_NOT), .b(EX461), .O(EX462) );
and2 gate( .a(N1476), .b(p186), .O(EX463) );
and2 gate( .a(N1504_NOT), .b(EX463), .O(EX464) );
and2 gate( .a(N1476_NOT), .b(p187), .O(EX465) );
and2 gate( .a(N1504), .b(EX465), .O(EX466) );
and2 gate( .a(N1476), .b(p188), .O(EX467) );
and2 gate( .a(N1504), .b(EX467), .O(EX468) );
or2  gate( .a(EX462), .b(EX464), .O(EX469) );
or2  gate( .a(EX466), .b(EX469), .O(EX470) );
or2  gate( .a(EX468), .b(EX470), .O(N1540) );
inv1 gate428( .a(N1513), .O(N1546) );
inv1 gate429( .a(N1521), .O(N1554) );
inv1 gate430( .a(N1526), .O(N1557) );
inv1 gate431( .a(N1520), .O(N1561) );
nand2 gate432( .a(N1484), .b(N1531), .O(N1567) );
inv1 gate( .a(N1481),.O(N1481_NOT) );
inv1 gate( .a(N1532),.O(N1532_NOT));
and2 gate( .a(N1481_NOT), .b(p189), .O(EX471) );
and2 gate( .a(N1532_NOT), .b(EX471), .O(EX472) );
and2 gate( .a(N1481), .b(p190), .O(EX473) );
and2 gate( .a(N1532_NOT), .b(EX473), .O(EX474) );
and2 gate( .a(N1481_NOT), .b(p191), .O(EX475) );
and2 gate( .a(N1532), .b(EX475), .O(EX476) );
and2 gate( .a(N1481), .b(p192), .O(EX477) );
and2 gate( .a(N1532), .b(EX477), .O(EX478) );
or2  gate( .a(EX472), .b(EX474), .O(EX479) );
or2  gate( .a(EX476), .b(EX479), .O(EX480) );
or2  gate( .a(EX478), .b(EX480), .O(N1568) );
inv1 gate434( .a(N1510), .O(N1569) );
inv1 gate435( .a(N1527), .O(N1571) );
inv1 gate436( .a(N1529), .O(N1576) );
buf1 gate437( .a(N1522), .O(N1588) );
inv1 gate438( .a(N1534), .O(N1591) );
inv1 gate439( .a(N1537), .O(N1593) );
nand2 gate440( .a(N1540), .b(N1530), .O(N1594) );
inv1 gate441( .a(N1540), .O(N1595) );
inv1 gate( .a(N1567),.O(N1567_NOT) );
inv1 gate( .a(N1568),.O(N1568_NOT));
and2 gate( .a(N1567_NOT), .b(p193), .O(EX481) );
and2 gate( .a(N1568_NOT), .b(EX481), .O(EX482) );
and2 gate( .a(N1567), .b(p194), .O(EX483) );
and2 gate( .a(N1568_NOT), .b(EX483), .O(EX484) );
and2 gate( .a(N1567_NOT), .b(p195), .O(EX485) );
and2 gate( .a(N1568), .b(EX485), .O(EX486) );
and2 gate( .a(N1567), .b(p196), .O(EX487) );
and2 gate( .a(N1568), .b(EX487), .O(EX488) );
or2  gate( .a(EX482), .b(EX484), .O(EX489) );
or2  gate( .a(EX486), .b(EX489), .O(EX490) );
or2  gate( .a(EX488), .b(EX490), .O(N1596) );
buf1 gate443( .a(N1517), .O(N1600) );
buf1 gate444( .a(N1517), .O(N1603) );
buf1 gate445( .a(N1522), .O(N1606) );
buf1 gate446( .a(N1522), .O(N1609) );
buf1 gate447( .a(N1514), .O(N1612) );
buf1 gate448( .a(N1514), .O(N1615) );
buf1 gate449( .a(N1557), .O(N1620) );
buf1 gate450( .a(N1554), .O(N1623) );
inv1 gate451( .a(N1571), .O(N1635) );
inv1 gate( .a(N1478),.O(N1478_NOT) );
inv1 gate( .a(N1595),.O(N1595_NOT));
and2 gate( .a(N1478_NOT), .b(p197), .O(EX491) );
and2 gate( .a(N1595_NOT), .b(EX491), .O(EX492) );
and2 gate( .a(N1478), .b(p198), .O(EX493) );
and2 gate( .a(N1595_NOT), .b(EX493), .O(EX494) );
and2 gate( .a(N1478_NOT), .b(p199), .O(EX495) );
and2 gate( .a(N1595), .b(EX495), .O(EX496) );
and2 gate( .a(N1478), .b(p200), .O(EX497) );
and2 gate( .a(N1595), .b(EX497), .O(EX498) );
or2  gate( .a(EX492), .b(EX494), .O(EX499) );
or2  gate( .a(EX496), .b(EX499), .O(EX500) );
or2  gate( .a(EX498), .b(EX500), .O(N1636) );
nand2 gate453( .a(N1576), .b(N1569), .O(N1638) );
inv1 gate454( .a(N1576), .O(N1639) );
buf1 gate455( .a(N1561), .O(N1640) );
buf1 gate456( .a(N1561), .O(N1643) );
buf1 gate457( .a(N1546), .O(N1647) );
buf1 gate458( .a(N1546), .O(N1651) );
buf1 gate459( .a(N1554), .O(N1658) );
buf1 gate460( .a(N1557), .O(N1661) );
buf1 gate461( .a(N1557), .O(N1664) );
nand2 gate462( .a(N1596), .b(N893), .O(N1671) );
inv1 gate463( .a(N1596), .O(N1672) );
inv1 gate464( .a(N1600), .O(N1675) );
inv1 gate465( .a(N1603), .O(N1677) );
nand2 gate466( .a(N1606), .b(N1217), .O(N1678) );
inv1 gate467( .a(N1606), .O(N1679) );
nand2 gate468( .a(N1609), .b(N1219), .O(N1680) );
inv1 gate469( .a(N1609), .O(N1681) );
inv1 gate470( .a(N1612), .O(N1682) );
inv1 gate471( .a(N1615), .O(N1683) );
inv1 gate( .a(N1594),.O(N1594_NOT) );
inv1 gate( .a(N1636),.O(N1636_NOT));
and2 gate( .a(N1594_NOT), .b(p201), .O(EX501) );
and2 gate( .a(N1636_NOT), .b(EX501), .O(EX502) );
and2 gate( .a(N1594), .b(p202), .O(EX503) );
and2 gate( .a(N1636_NOT), .b(EX503), .O(EX504) );
and2 gate( .a(N1594_NOT), .b(p203), .O(EX505) );
and2 gate( .a(N1636), .b(EX505), .O(EX506) );
and2 gate( .a(N1594), .b(p204), .O(EX507) );
and2 gate( .a(N1636), .b(EX507), .O(EX508) );
or2  gate( .a(EX502), .b(EX504), .O(EX509) );
or2  gate( .a(EX506), .b(EX509), .O(EX510) );
or2  gate( .a(EX508), .b(EX510), .O(N1685) );
inv1 gate( .a(N1510),.O(N1510_NOT) );
inv1 gate( .a(N1639),.O(N1639_NOT));
and2 gate( .a(N1510_NOT), .b(p205), .O(EX511) );
and2 gate( .a(N1639_NOT), .b(EX511), .O(EX512) );
and2 gate( .a(N1510), .b(p206), .O(EX513) );
and2 gate( .a(N1639_NOT), .b(EX513), .O(EX514) );
and2 gate( .a(N1510_NOT), .b(p207), .O(EX515) );
and2 gate( .a(N1639), .b(EX515), .O(EX516) );
and2 gate( .a(N1510), .b(p208), .O(EX517) );
and2 gate( .a(N1639), .b(EX517), .O(EX518) );
or2  gate( .a(EX512), .b(EX514), .O(EX519) );
or2  gate( .a(EX516), .b(EX519), .O(EX520) );
or2  gate( .a(EX518), .b(EX520), .O(N1688) );
buf1 gate474( .a(N1588), .O(N1697) );
buf1 gate475( .a(N1588), .O(N1701) );
nand2 gate476( .a(N643), .b(N1672), .O(N1706) );
inv1 gate477( .a(N1643), .O(N1707) );
inv1 gate( .a(N1647),.O(N1647_NOT) );
inv1 gate( .a(N1675),.O(N1675_NOT));
and2 gate( .a(N1647_NOT), .b(p209), .O(EX521) );
and2 gate( .a(N1675_NOT), .b(EX521), .O(EX522) );
and2 gate( .a(N1647), .b(p210), .O(EX523) );
and2 gate( .a(N1675_NOT), .b(EX523), .O(EX524) );
and2 gate( .a(N1647_NOT), .b(p211), .O(EX525) );
and2 gate( .a(N1675), .b(EX525), .O(EX526) );
and2 gate( .a(N1647), .b(p212), .O(EX527) );
and2 gate( .a(N1675), .b(EX527), .O(EX528) );
or2  gate( .a(EX522), .b(EX524), .O(EX529) );
or2  gate( .a(EX526), .b(EX529), .O(EX530) );
or2  gate( .a(EX528), .b(EX530), .O(N1708) );
inv1 gate479( .a(N1647), .O(N1709) );
nand2 gate480( .a(N1651), .b(N1677), .O(N1710) );
inv1 gate481( .a(N1651), .O(N1711) );
nand2 gate482( .a(N1028), .b(N1679), .O(N1712) );
inv1 gate( .a(N1031),.O(N1031_NOT) );
inv1 gate( .a(N1681),.O(N1681_NOT));
and2 gate( .a(N1031_NOT), .b(p213), .O(EX531) );
and2 gate( .a(N1681_NOT), .b(EX531), .O(EX532) );
and2 gate( .a(N1031), .b(p214), .O(EX533) );
and2 gate( .a(N1681_NOT), .b(EX533), .O(EX534) );
and2 gate( .a(N1031_NOT), .b(p215), .O(EX535) );
and2 gate( .a(N1681), .b(EX535), .O(EX536) );
and2 gate( .a(N1031), .b(p216), .O(EX537) );
and2 gate( .a(N1681), .b(EX537), .O(EX538) );
or2  gate( .a(EX532), .b(EX534), .O(EX539) );
or2  gate( .a(EX536), .b(EX539), .O(EX540) );
or2  gate( .a(EX538), .b(EX540), .O(N1713) );
buf1 gate484( .a(N1620), .O(N1714) );
buf1 gate485( .a(N1620), .O(N1717) );
inv1 gate( .a(N1658),.O(N1658_NOT) );
inv1 gate( .a(N1593),.O(N1593_NOT));
and2 gate( .a(N1658_NOT), .b(p217), .O(EX541) );
and2 gate( .a(N1593_NOT), .b(EX541), .O(EX542) );
and2 gate( .a(N1658), .b(p218), .O(EX543) );
and2 gate( .a(N1593_NOT), .b(EX543), .O(EX544) );
and2 gate( .a(N1658_NOT), .b(p219), .O(EX545) );
and2 gate( .a(N1593), .b(EX545), .O(EX546) );
and2 gate( .a(N1658), .b(p220), .O(EX547) );
and2 gate( .a(N1593), .b(EX547), .O(EX548) );
or2  gate( .a(EX542), .b(EX544), .O(EX549) );
or2  gate( .a(EX546), .b(EX549), .O(EX550) );
or2  gate( .a(EX548), .b(EX550), .O(N1720) );
inv1 gate487( .a(N1658), .O(N1721) );
inv1 gate( .a(N1638),.O(N1638_NOT) );
inv1 gate( .a(N1688),.O(N1688_NOT));
and2 gate( .a(N1638_NOT), .b(p221), .O(EX551) );
and2 gate( .a(N1688_NOT), .b(EX551), .O(EX552) );
and2 gate( .a(N1638), .b(p222), .O(EX553) );
and2 gate( .a(N1688_NOT), .b(EX553), .O(EX554) );
and2 gate( .a(N1638_NOT), .b(p223), .O(EX555) );
and2 gate( .a(N1688), .b(EX555), .O(EX556) );
and2 gate( .a(N1638), .b(p224), .O(EX557) );
and2 gate( .a(N1688), .b(EX557), .O(EX558) );
or2  gate( .a(EX552), .b(EX554), .O(EX559) );
or2  gate( .a(EX556), .b(EX559), .O(EX560) );
or2  gate( .a(EX558), .b(EX560), .O(N1723) );
inv1 gate489( .a(N1661), .O(N1727) );
inv1 gate490( .a(N1640), .O(N1728) );
inv1 gate491( .a(N1664), .O(N1730) );
buf1 gate492( .a(N1623), .O(N1731) );
buf1 gate493( .a(N1623), .O(N1734) );
inv1 gate( .a(N1685),.O(N1685_NOT) );
inv1 gate( .a(N1528),.O(N1528_NOT));
and2 gate( .a(N1685_NOT), .b(p225), .O(EX561) );
and2 gate( .a(N1528_NOT), .b(EX561), .O(EX562) );
and2 gate( .a(N1685), .b(p226), .O(EX563) );
and2 gate( .a(N1528_NOT), .b(EX563), .O(EX564) );
and2 gate( .a(N1685_NOT), .b(p227), .O(EX565) );
and2 gate( .a(N1528), .b(EX565), .O(EX566) );
and2 gate( .a(N1685), .b(p228), .O(EX567) );
and2 gate( .a(N1528), .b(EX567), .O(EX568) );
or2  gate( .a(EX562), .b(EX564), .O(EX569) );
or2  gate( .a(EX566), .b(EX569), .O(EX570) );
or2  gate( .a(EX568), .b(EX570), .O(N1740) );
inv1 gate495( .a(N1685), .O(N1741) );
nand2 gate496( .a(N1671), .b(N1706), .O(N1742) );
inv1 gate( .a(N1600),.O(N1600_NOT) );
inv1 gate( .a(N1709),.O(N1709_NOT));
and2 gate( .a(N1600_NOT), .b(p229), .O(EX571) );
and2 gate( .a(N1709_NOT), .b(EX571), .O(EX572) );
and2 gate( .a(N1600), .b(p230), .O(EX573) );
and2 gate( .a(N1709_NOT), .b(EX573), .O(EX574) );
and2 gate( .a(N1600_NOT), .b(p231), .O(EX575) );
and2 gate( .a(N1709), .b(EX575), .O(EX576) );
and2 gate( .a(N1600), .b(p232), .O(EX577) );
and2 gate( .a(N1709), .b(EX577), .O(EX578) );
or2  gate( .a(EX572), .b(EX574), .O(EX579) );
or2  gate( .a(EX576), .b(EX579), .O(EX580) );
or2  gate( .a(EX578), .b(EX580), .O(N1746) );
nand2 gate498( .a(N1603), .b(N1711), .O(N1747) );
inv1 gate( .a(N1678),.O(N1678_NOT) );
inv1 gate( .a(N1712),.O(N1712_NOT));
and2 gate( .a(N1678_NOT), .b(p233), .O(EX581) );
and2 gate( .a(N1712_NOT), .b(EX581), .O(EX582) );
and2 gate( .a(N1678), .b(p234), .O(EX583) );
and2 gate( .a(N1712_NOT), .b(EX583), .O(EX584) );
and2 gate( .a(N1678_NOT), .b(p235), .O(EX585) );
and2 gate( .a(N1712), .b(EX585), .O(EX586) );
and2 gate( .a(N1678), .b(p236), .O(EX587) );
and2 gate( .a(N1712), .b(EX587), .O(EX588) );
or2  gate( .a(EX582), .b(EX584), .O(EX589) );
or2  gate( .a(EX586), .b(EX589), .O(EX590) );
or2  gate( .a(EX588), .b(EX590), .O(N1748) );
nand2 gate500( .a(N1680), .b(N1713), .O(N1751) );
inv1 gate( .a(N1537),.O(N1537_NOT) );
inv1 gate( .a(N1721),.O(N1721_NOT));
and2 gate( .a(N1537_NOT), .b(p237), .O(EX591) );
and2 gate( .a(N1721_NOT), .b(EX591), .O(EX592) );
and2 gate( .a(N1537), .b(p238), .O(EX593) );
and2 gate( .a(N1721_NOT), .b(EX593), .O(EX594) );
and2 gate( .a(N1537_NOT), .b(p239), .O(EX595) );
and2 gate( .a(N1721), .b(EX595), .O(EX596) );
and2 gate( .a(N1537), .b(p240), .O(EX597) );
and2 gate( .a(N1721), .b(EX597), .O(EX598) );
or2  gate( .a(EX592), .b(EX594), .O(EX599) );
or2  gate( .a(EX596), .b(EX599), .O(EX600) );
or2  gate( .a(EX598), .b(EX600), .O(N1759) );
inv1 gate502( .a(N1697), .O(N1761) );
inv1 gate( .a(N1697),.O(N1697_NOT) );
inv1 gate( .a(N1727),.O(N1727_NOT));
and2 gate( .a(N1697_NOT), .b(p241), .O(EX601) );
and2 gate( .a(N1727_NOT), .b(EX601), .O(EX602) );
and2 gate( .a(N1697), .b(p242), .O(EX603) );
and2 gate( .a(N1727_NOT), .b(EX603), .O(EX604) );
and2 gate( .a(N1697_NOT), .b(p243), .O(EX605) );
and2 gate( .a(N1727), .b(EX605), .O(EX606) );
and2 gate( .a(N1697), .b(p244), .O(EX607) );
and2 gate( .a(N1727), .b(EX607), .O(EX608) );
or2  gate( .a(EX602), .b(EX604), .O(EX609) );
or2  gate( .a(EX606), .b(EX609), .O(EX610) );
or2  gate( .a(EX608), .b(EX610), .O(N1762) );
inv1 gate504( .a(N1701), .O(N1763) );
nand2 gate505( .a(N1701), .b(N1730), .O(N1764) );
inv1 gate506( .a(N1717), .O(N1768) );
nand2 gate507( .a(N1472), .b(N1741), .O(N1769) );
nand2 gate508( .a(N1723), .b(N1413), .O(N1772) );
inv1 gate509( .a(N1723), .O(N1773) );
inv1 gate( .a(N1708),.O(N1708_NOT) );
inv1 gate( .a(N1746),.O(N1746_NOT));
and2 gate( .a(N1708_NOT), .b(p245), .O(EX611) );
and2 gate( .a(N1746_NOT), .b(EX611), .O(EX612) );
and2 gate( .a(N1708), .b(p246), .O(EX613) );
and2 gate( .a(N1746_NOT), .b(EX613), .O(EX614) );
and2 gate( .a(N1708_NOT), .b(p247), .O(EX615) );
and2 gate( .a(N1746), .b(EX615), .O(EX616) );
and2 gate( .a(N1708), .b(p248), .O(EX617) );
and2 gate( .a(N1746), .b(EX617), .O(EX618) );
or2  gate( .a(EX612), .b(EX614), .O(EX619) );
or2  gate( .a(EX616), .b(EX619), .O(EX620) );
or2  gate( .a(EX618), .b(EX620), .O(N1774) );
nand2 gate511( .a(N1710), .b(N1747), .O(N1777) );
inv1 gate512( .a(N1731), .O(N1783) );
nand2 gate513( .a(N1731), .b(N1682), .O(N1784) );
inv1 gate514( .a(N1714), .O(N1785) );
inv1 gate515( .a(N1734), .O(N1786) );
nand2 gate516( .a(N1734), .b(N1683), .O(N1787) );
nand2 gate517( .a(N1720), .b(N1759), .O(N1788) );
nand2 gate518( .a(N1661), .b(N1761), .O(N1791) );
inv1 gate( .a(N1664),.O(N1664_NOT) );
inv1 gate( .a(N1763),.O(N1763_NOT));
and2 gate( .a(N1664_NOT), .b(p249), .O(EX621) );
and2 gate( .a(N1763_NOT), .b(EX621), .O(EX622) );
and2 gate( .a(N1664), .b(p250), .O(EX623) );
and2 gate( .a(N1763_NOT), .b(EX623), .O(EX624) );
and2 gate( .a(N1664_NOT), .b(p251), .O(EX625) );
and2 gate( .a(N1763), .b(EX625), .O(EX626) );
and2 gate( .a(N1664), .b(p252), .O(EX627) );
and2 gate( .a(N1763), .b(EX627), .O(EX628) );
or2  gate( .a(EX622), .b(EX624), .O(EX629) );
or2  gate( .a(EX626), .b(EX629), .O(EX630) );
or2  gate( .a(EX628), .b(EX630), .O(N1792) );
nand2 gate520( .a(N1751), .b(N1155), .O(N1795) );
inv1 gate521( .a(N1751), .O(N1796) );
nand2 gate522( .a(N1740), .b(N1769), .O(N1798) );
inv1 gate( .a(N1334),.O(N1334_NOT) );
inv1 gate( .a(N1773),.O(N1773_NOT));
and2 gate( .a(N1334_NOT), .b(p253), .O(EX631) );
and2 gate( .a(N1773_NOT), .b(EX631), .O(EX632) );
and2 gate( .a(N1334), .b(p254), .O(EX633) );
and2 gate( .a(N1773_NOT), .b(EX633), .O(EX634) );
and2 gate( .a(N1334_NOT), .b(p255), .O(EX635) );
and2 gate( .a(N1773), .b(EX635), .O(EX636) );
and2 gate( .a(N1334), .b(p256), .O(EX637) );
and2 gate( .a(N1773), .b(EX637), .O(EX638) );
or2  gate( .a(EX632), .b(EX634), .O(EX639) );
or2  gate( .a(EX636), .b(EX639), .O(EX640) );
or2  gate( .a(EX638), .b(EX640), .O(N1801) );
nand2 gate524( .a(N1742), .b(N290), .O(N1802) );
inv1 gate525( .a(N1748), .O(N1807) );
nand2 gate526( .a(N1748), .b(N1218), .O(N1808) );
nand2 gate527( .a(N1612), .b(N1783), .O(N1809) );
nand2 gate528( .a(N1615), .b(N1786), .O(N1810) );
nand2 gate529( .a(N1791), .b(N1762), .O(N1812) );
nand2 gate530( .a(N1792), .b(N1764), .O(N1815) );
buf1 gate531( .a(N1742), .O(N1818) );
inv1 gate( .a(N1777),.O(N1777_NOT) );
inv1 gate( .a(N1490),.O(N1490_NOT));
and2 gate( .a(N1777_NOT), .b(p257), .O(EX641) );
and2 gate( .a(N1490_NOT), .b(EX641), .O(EX642) );
and2 gate( .a(N1777), .b(p258), .O(EX643) );
and2 gate( .a(N1490_NOT), .b(EX643), .O(EX644) );
and2 gate( .a(N1777_NOT), .b(p259), .O(EX645) );
and2 gate( .a(N1490), .b(EX645), .O(EX646) );
and2 gate( .a(N1777), .b(p260), .O(EX647) );
and2 gate( .a(N1490), .b(EX647), .O(EX648) );
or2  gate( .a(EX642), .b(EX644), .O(EX649) );
or2  gate( .a(EX646), .b(EX649), .O(EX650) );
or2  gate( .a(EX648), .b(EX650), .O(N1821) );
inv1 gate533( .a(N1777), .O(N1822) );
nand2 gate534( .a(N1774), .b(N1491), .O(N1823) );
inv1 gate535( .a(N1774), .O(N1824) );
nand2 gate536( .a(N962), .b(N1796), .O(N1825) );
nand2 gate537( .a(N1788), .b(N1409), .O(N1826) );
inv1 gate538( .a(N1788), .O(N1827) );
nand2 gate539( .a(N1772), .b(N1801), .O(N1830) );
nand2 gate540( .a(N959), .b(N1807), .O(N1837) );
nand2 gate541( .a(N1809), .b(N1784), .O(N1838) );
nand2 gate542( .a(N1810), .b(N1787), .O(N1841) );
nand2 gate543( .a(N1419), .b(N1822), .O(N1848) );
nand2 gate544( .a(N1416), .b(N1824), .O(N1849) );
nand2 gate545( .a(N1795), .b(N1825), .O(N1850) );
nand2 gate546( .a(N1319), .b(N1827), .O(N1852) );
inv1 gate( .a(N1815),.O(N1815_NOT) );
inv1 gate( .a(N1707),.O(N1707_NOT));
and2 gate( .a(N1815_NOT), .b(p261), .O(EX651) );
and2 gate( .a(N1707_NOT), .b(EX651), .O(EX652) );
and2 gate( .a(N1815), .b(p262), .O(EX653) );
and2 gate( .a(N1707_NOT), .b(EX653), .O(EX654) );
and2 gate( .a(N1815_NOT), .b(p263), .O(EX655) );
and2 gate( .a(N1707), .b(EX655), .O(EX656) );
and2 gate( .a(N1815), .b(p264), .O(EX657) );
and2 gate( .a(N1707), .b(EX657), .O(EX658) );
or2  gate( .a(EX652), .b(EX654), .O(EX659) );
or2  gate( .a(EX656), .b(EX659), .O(EX660) );
or2  gate( .a(EX658), .b(EX660), .O(N1855) );
inv1 gate548( .a(N1815), .O(N1856) );
inv1 gate549( .a(N1818), .O(N1857) );
nand2 gate550( .a(N1798), .b(N290), .O(N1858) );
inv1 gate551( .a(N1812), .O(N1864) );
nand2 gate552( .a(N1812), .b(N1728), .O(N1865) );
buf1 gate553( .a(N1798), .O(N1866) );
buf1 gate554( .a(N1802), .O(N1869) );
buf1 gate555( .a(N1802), .O(N1872) );
nand2 gate556( .a(N1808), .b(N1837), .O(N1875) );
nand2 gate557( .a(N1821), .b(N1848), .O(N1878) );
nand2 gate558( .a(N1823), .b(N1849), .O(N1879) );
nand2 gate559( .a(N1841), .b(N1768), .O(N1882) );
inv1 gate560( .a(N1841), .O(N1883) );
nand2 gate561( .a(N1826), .b(N1852), .O(N1884) );
nand2 gate562( .a(N1643), .b(N1856), .O(N1885) );
nand2 gate563( .a(N1830), .b(N290), .O(N1889) );
inv1 gate564( .a(N1838), .O(N1895) );
nand2 gate565( .a(N1838), .b(N1785), .O(N1896) );
nand2 gate566( .a(N1640), .b(N1864), .O(N1897) );
inv1 gate567( .a(N1850), .O(N1898) );
buf1 gate568( .a(N1830), .O(N1902) );
inv1 gate569( .a(N1878), .O(N1910) );
nand2 gate570( .a(N1717), .b(N1883), .O(N1911) );
inv1 gate571( .a(N1884), .O(N1912) );
inv1 gate( .a(N1855),.O(N1855_NOT) );
inv1 gate( .a(N1885),.O(N1885_NOT));
and2 gate( .a(N1855_NOT), .b(p265), .O(EX661) );
and2 gate( .a(N1885_NOT), .b(EX661), .O(EX662) );
and2 gate( .a(N1855), .b(p266), .O(EX663) );
and2 gate( .a(N1885_NOT), .b(EX663), .O(EX664) );
and2 gate( .a(N1855_NOT), .b(p267), .O(EX665) );
and2 gate( .a(N1885), .b(EX665), .O(EX666) );
and2 gate( .a(N1855), .b(p268), .O(EX667) );
and2 gate( .a(N1885), .b(EX667), .O(EX668) );
or2  gate( .a(EX662), .b(EX664), .O(EX669) );
or2  gate( .a(EX666), .b(EX669), .O(EX670) );
or2  gate( .a(EX668), .b(EX670), .O(N1913) );
inv1 gate573( .a(N1866), .O(N1915) );
nand2 gate574( .a(N1872), .b(N919), .O(N1919) );
inv1 gate575( .a(N1872), .O(N1920) );
nand2 gate576( .a(N1869), .b(N920), .O(N1921) );
inv1 gate577( .a(N1869), .O(N1922) );
inv1 gate578( .a(N1875), .O(N1923) );
nand2 gate579( .a(N1714), .b(N1895), .O(N1924) );
buf1 gate580( .a(N1858), .O(N1927) );
buf1 gate581( .a(N1858), .O(N1930) );
nand2 gate582( .a(N1865), .b(N1897), .O(N1933) );
nand2 gate583( .a(N1882), .b(N1911), .O(N1936) );
inv1 gate584( .a(N1898), .O(N1937) );
inv1 gate585( .a(N1902), .O(N1938) );
inv1 gate( .a(N679),.O(N679_NOT) );
inv1 gate( .a(N1920),.O(N1920_NOT));
and2 gate( .a(N679_NOT), .b(p269), .O(EX671) );
and2 gate( .a(N1920_NOT), .b(EX671), .O(EX672) );
and2 gate( .a(N679), .b(p270), .O(EX673) );
and2 gate( .a(N1920_NOT), .b(EX673), .O(EX674) );
and2 gate( .a(N679_NOT), .b(p271), .O(EX675) );
and2 gate( .a(N1920), .b(EX675), .O(EX676) );
and2 gate( .a(N679), .b(p272), .O(EX677) );
and2 gate( .a(N1920), .b(EX677), .O(EX678) );
or2  gate( .a(EX672), .b(EX674), .O(EX679) );
or2  gate( .a(EX676), .b(EX679), .O(EX680) );
or2  gate( .a(EX678), .b(EX680), .O(N1941) );
inv1 gate( .a(N676),.O(N676_NOT) );
inv1 gate( .a(N1922),.O(N1922_NOT));
and2 gate( .a(N676_NOT), .b(p273), .O(EX681) );
and2 gate( .a(N1922_NOT), .b(EX681), .O(EX682) );
and2 gate( .a(N676), .b(p274), .O(EX683) );
and2 gate( .a(N1922_NOT), .b(EX683), .O(EX684) );
and2 gate( .a(N676_NOT), .b(p275), .O(EX685) );
and2 gate( .a(N1922), .b(EX685), .O(EX686) );
and2 gate( .a(N676), .b(p276), .O(EX687) );
and2 gate( .a(N1922), .b(EX687), .O(EX688) );
or2  gate( .a(EX682), .b(EX684), .O(EX689) );
or2  gate( .a(EX686), .b(EX689), .O(EX690) );
or2  gate( .a(EX688), .b(EX690), .O(N1942) );
buf1 gate588( .a(N1879), .O(N1944) );
inv1 gate589( .a(N1913), .O(N1947) );
buf1 gate590( .a(N1889), .O(N1950) );
buf1 gate591( .a(N1889), .O(N1953) );
buf1 gate592( .a(N1879), .O(N1958) );
nand2 gate593( .a(N1896), .b(N1924), .O(N1961) );
and2 gate594( .a(N1910), .b(N601), .O(N1965) );
and2 gate595( .a(N602), .b(N1912), .O(N1968) );
nand2 gate596( .a(N1930), .b(N917), .O(N1975) );
inv1 gate597( .a(N1930), .O(N1976) );
nand2 gate598( .a(N1927), .b(N918), .O(N1977) );
inv1 gate599( .a(N1927), .O(N1978) );
nand2 gate600( .a(N1919), .b(N1941), .O(N1979) );
inv1 gate( .a(N1921),.O(N1921_NOT) );
inv1 gate( .a(N1942),.O(N1942_NOT));
and2 gate( .a(N1921_NOT), .b(p277), .O(EX691) );
and2 gate( .a(N1942_NOT), .b(EX691), .O(EX692) );
and2 gate( .a(N1921), .b(p278), .O(EX693) );
and2 gate( .a(N1942_NOT), .b(EX693), .O(EX694) );
and2 gate( .a(N1921_NOT), .b(p279), .O(EX695) );
and2 gate( .a(N1942), .b(EX695), .O(EX696) );
and2 gate( .a(N1921), .b(p280), .O(EX697) );
and2 gate( .a(N1942), .b(EX697), .O(EX698) );
or2  gate( .a(EX692), .b(EX694), .O(EX699) );
or2  gate( .a(EX696), .b(EX699), .O(EX700) );
or2  gate( .a(EX698), .b(EX700), .O(N1980) );
inv1 gate602( .a(N1933), .O(N1985) );
inv1 gate603( .a(N1936), .O(N1987) );
inv1 gate604( .a(N1944), .O(N1999) );
nand2 gate605( .a(N1944), .b(N1937), .O(N2000) );
inv1 gate606( .a(N1947), .O(N2002) );
inv1 gate( .a(N1947),.O(N1947_NOT) );
inv1 gate( .a(N1499),.O(N1499_NOT));
and2 gate( .a(N1947_NOT), .b(p281), .O(EX701) );
and2 gate( .a(N1499_NOT), .b(EX701), .O(EX702) );
and2 gate( .a(N1947), .b(p282), .O(EX703) );
and2 gate( .a(N1499_NOT), .b(EX703), .O(EX704) );
and2 gate( .a(N1947_NOT), .b(p283), .O(EX705) );
and2 gate( .a(N1499), .b(EX705), .O(EX706) );
and2 gate( .a(N1947), .b(p284), .O(EX707) );
and2 gate( .a(N1499), .b(EX707), .O(EX708) );
or2  gate( .a(EX702), .b(EX704), .O(EX709) );
or2  gate( .a(EX706), .b(EX709), .O(EX710) );
or2  gate( .a(EX708), .b(EX710), .O(N2003) );
nand2 gate608( .a(N1953), .b(N1350), .O(N2004) );
inv1 gate609( .a(N1953), .O(N2005) );
nand2 gate610( .a(N1950), .b(N1351), .O(N2006) );
inv1 gate611( .a(N1950), .O(N2007) );
inv1 gate( .a(N673),.O(N673_NOT) );
inv1 gate( .a(N1976),.O(N1976_NOT));
and2 gate( .a(N673_NOT), .b(p285), .O(EX711) );
and2 gate( .a(N1976_NOT), .b(EX711), .O(EX712) );
and2 gate( .a(N673), .b(p286), .O(EX713) );
and2 gate( .a(N1976_NOT), .b(EX713), .O(EX714) );
and2 gate( .a(N673_NOT), .b(p287), .O(EX715) );
and2 gate( .a(N1976), .b(EX715), .O(EX716) );
and2 gate( .a(N673), .b(p288), .O(EX717) );
and2 gate( .a(N1976), .b(EX717), .O(EX718) );
or2  gate( .a(EX712), .b(EX714), .O(EX719) );
or2  gate( .a(EX716), .b(EX719), .O(EX720) );
or2  gate( .a(EX718), .b(EX720), .O(N2008) );
nand2 gate613( .a(N670), .b(N1978), .O(N2009) );
inv1 gate614( .a(N1979), .O(N2012) );
inv1 gate615( .a(N1958), .O(N2013) );
nand2 gate616( .a(N1958), .b(N1923), .O(N2014) );
inv1 gate617( .a(N1961), .O(N2015) );
nand2 gate618( .a(N1961), .b(N1635), .O(N2016) );
inv1 gate619( .a(N1965), .O(N2018) );
inv1 gate620( .a(N1968), .O(N2019) );
nand2 gate621( .a(N1898), .b(N1999), .O(N2020) );
inv1 gate622( .a(N1987), .O(N2021) );
nand2 gate623( .a(N1987), .b(N1591), .O(N2022) );
nand2 gate624( .a(N1440), .b(N2002), .O(N2023) );
nand2 gate625( .a(N1261), .b(N2005), .O(N2024) );
inv1 gate( .a(N1258),.O(N1258_NOT) );
inv1 gate( .a(N2007),.O(N2007_NOT));
and2 gate( .a(N1258_NOT), .b(p289), .O(EX721) );
and2 gate( .a(N2007_NOT), .b(EX721), .O(EX722) );
and2 gate( .a(N1258), .b(p290), .O(EX723) );
and2 gate( .a(N2007_NOT), .b(EX723), .O(EX724) );
and2 gate( .a(N1258_NOT), .b(p291), .O(EX725) );
and2 gate( .a(N2007), .b(EX725), .O(EX726) );
and2 gate( .a(N1258), .b(p292), .O(EX727) );
and2 gate( .a(N2007), .b(EX727), .O(EX728) );
or2  gate( .a(EX722), .b(EX724), .O(EX729) );
or2  gate( .a(EX726), .b(EX729), .O(EX730) );
or2  gate( .a(EX728), .b(EX730), .O(N2025) );
nand2 gate627( .a(N1975), .b(N2008), .O(N2026) );
inv1 gate( .a(N1977),.O(N1977_NOT) );
inv1 gate( .a(N2009),.O(N2009_NOT));
and2 gate( .a(N1977_NOT), .b(p293), .O(EX731) );
and2 gate( .a(N2009_NOT), .b(EX731), .O(EX732) );
and2 gate( .a(N1977), .b(p294), .O(EX733) );
and2 gate( .a(N2009_NOT), .b(EX733), .O(EX734) );
and2 gate( .a(N1977_NOT), .b(p295), .O(EX735) );
and2 gate( .a(N2009), .b(EX735), .O(EX736) );
and2 gate( .a(N1977), .b(p296), .O(EX737) );
and2 gate( .a(N2009), .b(EX737), .O(EX738) );
or2  gate( .a(EX732), .b(EX734), .O(EX739) );
or2  gate( .a(EX736), .b(EX739), .O(EX740) );
or2  gate( .a(EX738), .b(EX740), .O(N2027) );
inv1 gate629( .a(N1980), .O(N2030) );
buf1 gate630( .a(N1980), .O(N2033) );
nand2 gate631( .a(N1875), .b(N2013), .O(N2036) );
nand2 gate632( .a(N1571), .b(N2015), .O(N2037) );
nand2 gate633( .a(N2020), .b(N2000), .O(N2038) );
inv1 gate( .a(N1534),.O(N1534_NOT) );
inv1 gate( .a(N2021),.O(N2021_NOT));
and2 gate( .a(N1534_NOT), .b(p297), .O(EX741) );
and2 gate( .a(N2021_NOT), .b(EX741), .O(EX742) );
and2 gate( .a(N1534), .b(p298), .O(EX743) );
and2 gate( .a(N2021_NOT), .b(EX743), .O(EX744) );
and2 gate( .a(N1534_NOT), .b(p299), .O(EX745) );
and2 gate( .a(N2021), .b(EX745), .O(EX746) );
and2 gate( .a(N1534), .b(p300), .O(EX747) );
and2 gate( .a(N2021), .b(EX747), .O(EX748) );
or2  gate( .a(EX742), .b(EX744), .O(EX749) );
or2  gate( .a(EX746), .b(EX749), .O(EX750) );
or2  gate( .a(EX748), .b(EX750), .O(N2039) );
nand2 gate635( .a(N2023), .b(N2003), .O(N2040) );
inv1 gate( .a(N2004),.O(N2004_NOT) );
inv1 gate( .a(N2024),.O(N2024_NOT));
and2 gate( .a(N2004_NOT), .b(p301), .O(EX751) );
and2 gate( .a(N2024_NOT), .b(EX751), .O(EX752) );
and2 gate( .a(N2004), .b(p302), .O(EX753) );
and2 gate( .a(N2024_NOT), .b(EX753), .O(EX754) );
and2 gate( .a(N2004_NOT), .b(p303), .O(EX755) );
and2 gate( .a(N2024), .b(EX755), .O(EX756) );
and2 gate( .a(N2004), .b(p304), .O(EX757) );
and2 gate( .a(N2024), .b(EX757), .O(EX758) );
or2  gate( .a(EX752), .b(EX754), .O(EX759) );
or2  gate( .a(EX756), .b(EX759), .O(EX760) );
or2  gate( .a(EX758), .b(EX760), .O(N2041) );
nand2 gate637( .a(N2006), .b(N2025), .O(N2042) );
inv1 gate638( .a(N2026), .O(N2047) );
nand2 gate639( .a(N2036), .b(N2014), .O(N2052) );
nand2 gate640( .a(N2037), .b(N2016), .O(N2055) );
inv1 gate641( .a(N2038), .O(N2060) );
nand2 gate642( .a(N2039), .b(N2022), .O(N2061) );
nand2 gate643( .a(N2040), .b(N290), .O(N2062) );
inv1 gate644( .a(N2041), .O(N2067) );
inv1 gate645( .a(N2027), .O(N2068) );
buf1 gate646( .a(N2027), .O(N2071) );
inv1 gate647( .a(N2052), .O(N2076) );
inv1 gate648( .a(N2055), .O(N2077) );
inv1 gate( .a(N2060),.O(N2060_NOT) );
inv1 gate( .a(N290),.O(N290_NOT));
and2 gate( .a(N2060_NOT), .b(p305), .O(EX761) );
and2 gate( .a(N290_NOT), .b(EX761), .O(EX762) );
and2 gate( .a(N2060), .b(p306), .O(EX763) );
and2 gate( .a(N290_NOT), .b(EX763), .O(EX764) );
and2 gate( .a(N2060_NOT), .b(p307), .O(EX765) );
and2 gate( .a(N290), .b(EX765), .O(EX766) );
and2 gate( .a(N2060), .b(p308), .O(EX767) );
and2 gate( .a(N290), .b(EX767), .O(EX768) );
or2  gate( .a(EX762), .b(EX764), .O(EX769) );
or2  gate( .a(EX766), .b(EX769), .O(EX770) );
or2  gate( .a(EX768), .b(EX770), .O(N2078) );
nand2 gate650( .a(N2061), .b(N290), .O(N2081) );
inv1 gate651( .a(N2042), .O(N2086) );
buf1 gate652( .a(N2042), .O(N2089) );
and2 gate653( .a(N2030), .b(N2068), .O(N2104) );
and2 gate654( .a(N2033), .b(N2068), .O(N2119) );
and2 gate655( .a(N2030), .b(N2071), .O(N2129) );
and2 gate656( .a(N2033), .b(N2071), .O(N2143) );
buf1 gate657( .a(N2062), .O(N2148) );
buf1 gate658( .a(N2062), .O(N2151) );
buf1 gate659( .a(N2078), .O(N2196) );
buf1 gate660( .a(N2078), .O(N2199) );
buf1 gate661( .a(N2081), .O(N2202) );
buf1 gate662( .a(N2081), .O(N2205) );
nand2 gate663( .a(N2151), .b(N915), .O(N2214) );
inv1 gate664( .a(N2151), .O(N2215) );
nand2 gate665( .a(N2148), .b(N916), .O(N2216) );
inv1 gate666( .a(N2148), .O(N2217) );
inv1 gate( .a(N2199),.O(N2199_NOT) );
inv1 gate( .a(N1348),.O(N1348_NOT));
and2 gate( .a(N2199_NOT), .b(p309), .O(EX771) );
and2 gate( .a(N1348_NOT), .b(EX771), .O(EX772) );
and2 gate( .a(N2199), .b(p310), .O(EX773) );
and2 gate( .a(N1348_NOT), .b(EX773), .O(EX774) );
and2 gate( .a(N2199_NOT), .b(p311), .O(EX775) );
and2 gate( .a(N1348), .b(EX775), .O(EX776) );
and2 gate( .a(N2199), .b(p312), .O(EX777) );
and2 gate( .a(N1348), .b(EX777), .O(EX778) );
or2  gate( .a(EX772), .b(EX774), .O(EX779) );
or2  gate( .a(EX776), .b(EX779), .O(EX780) );
or2  gate( .a(EX778), .b(EX780), .O(N2222) );
inv1 gate668( .a(N2199), .O(N2223) );
inv1 gate( .a(N2196),.O(N2196_NOT) );
inv1 gate( .a(N1349),.O(N1349_NOT));
and2 gate( .a(N2196_NOT), .b(p313), .O(EX781) );
and2 gate( .a(N1349_NOT), .b(EX781), .O(EX782) );
and2 gate( .a(N2196), .b(p314), .O(EX783) );
and2 gate( .a(N1349_NOT), .b(EX783), .O(EX784) );
and2 gate( .a(N2196_NOT), .b(p315), .O(EX785) );
and2 gate( .a(N1349), .b(EX785), .O(EX786) );
and2 gate( .a(N2196), .b(p316), .O(EX787) );
and2 gate( .a(N1349), .b(EX787), .O(EX788) );
or2  gate( .a(EX782), .b(EX784), .O(EX789) );
or2  gate( .a(EX786), .b(EX789), .O(EX790) );
or2  gate( .a(EX788), .b(EX790), .O(N2224) );
inv1 gate670( .a(N2196), .O(N2225) );
nand2 gate671( .a(N2205), .b(N913), .O(N2226) );
inv1 gate672( .a(N2205), .O(N2227) );
nand2 gate673( .a(N2202), .b(N914), .O(N2228) );
inv1 gate674( .a(N2202), .O(N2229) );
inv1 gate( .a(N667),.O(N667_NOT) );
inv1 gate( .a(N2215),.O(N2215_NOT));
and2 gate( .a(N667_NOT), .b(p317), .O(EX791) );
and2 gate( .a(N2215_NOT), .b(EX791), .O(EX792) );
and2 gate( .a(N667), .b(p318), .O(EX793) );
and2 gate( .a(N2215_NOT), .b(EX793), .O(EX794) );
and2 gate( .a(N667_NOT), .b(p319), .O(EX795) );
and2 gate( .a(N2215), .b(EX795), .O(EX796) );
and2 gate( .a(N667), .b(p320), .O(EX797) );
and2 gate( .a(N2215), .b(EX797), .O(EX798) );
or2  gate( .a(EX792), .b(EX794), .O(EX799) );
or2  gate( .a(EX796), .b(EX799), .O(EX800) );
or2  gate( .a(EX798), .b(EX800), .O(N2230) );
inv1 gate( .a(N664),.O(N664_NOT) );
inv1 gate( .a(N2217),.O(N2217_NOT));
and2 gate( .a(N664_NOT), .b(p321), .O(EX801) );
and2 gate( .a(N2217_NOT), .b(EX801), .O(EX802) );
and2 gate( .a(N664), .b(p322), .O(EX803) );
and2 gate( .a(N2217_NOT), .b(EX803), .O(EX804) );
and2 gate( .a(N664_NOT), .b(p323), .O(EX805) );
and2 gate( .a(N2217), .b(EX805), .O(EX806) );
and2 gate( .a(N664), .b(p324), .O(EX807) );
and2 gate( .a(N2217), .b(EX807), .O(EX808) );
or2  gate( .a(EX802), .b(EX804), .O(EX809) );
or2  gate( .a(EX806), .b(EX809), .O(EX810) );
or2  gate( .a(EX808), .b(EX810), .O(N2231) );
inv1 gate( .a(N1255),.O(N1255_NOT) );
inv1 gate( .a(N2223),.O(N2223_NOT));
and2 gate( .a(N1255_NOT), .b(p325), .O(EX811) );
and2 gate( .a(N2223_NOT), .b(EX811), .O(EX812) );
and2 gate( .a(N1255), .b(p326), .O(EX813) );
and2 gate( .a(N2223_NOT), .b(EX813), .O(EX814) );
and2 gate( .a(N1255_NOT), .b(p327), .O(EX815) );
and2 gate( .a(N2223), .b(EX815), .O(EX816) );
and2 gate( .a(N1255), .b(p328), .O(EX817) );
and2 gate( .a(N2223), .b(EX817), .O(EX818) );
or2  gate( .a(EX812), .b(EX814), .O(EX819) );
or2  gate( .a(EX816), .b(EX819), .O(EX820) );
or2  gate( .a(EX818), .b(EX820), .O(N2232) );
inv1 gate( .a(N1252),.O(N1252_NOT) );
inv1 gate( .a(N2225),.O(N2225_NOT));
and2 gate( .a(N1252_NOT), .b(p329), .O(EX821) );
and2 gate( .a(N2225_NOT), .b(EX821), .O(EX822) );
and2 gate( .a(N1252), .b(p330), .O(EX823) );
and2 gate( .a(N2225_NOT), .b(EX823), .O(EX824) );
and2 gate( .a(N1252_NOT), .b(p331), .O(EX825) );
and2 gate( .a(N2225), .b(EX825), .O(EX826) );
and2 gate( .a(N1252), .b(p332), .O(EX827) );
and2 gate( .a(N2225), .b(EX827), .O(EX828) );
or2  gate( .a(EX822), .b(EX824), .O(EX829) );
or2  gate( .a(EX826), .b(EX829), .O(EX830) );
or2  gate( .a(EX828), .b(EX830), .O(N2233) );
nand2 gate679( .a(N661), .b(N2227), .O(N2234) );
nand2 gate680( .a(N658), .b(N2229), .O(N2235) );
nand2 gate681( .a(N2214), .b(N2230), .O(N2236) );
nand2 gate682( .a(N2216), .b(N2231), .O(N2237) );
nand2 gate683( .a(N2222), .b(N2232), .O(N2240) );
nand2 gate684( .a(N2224), .b(N2233), .O(N2241) );
nand2 gate685( .a(N2226), .b(N2234), .O(N2244) );
inv1 gate( .a(N2228),.O(N2228_NOT) );
inv1 gate( .a(N2235),.O(N2235_NOT));
and2 gate( .a(N2228_NOT), .b(p333), .O(EX831) );
and2 gate( .a(N2235_NOT), .b(EX831), .O(EX832) );
and2 gate( .a(N2228), .b(p334), .O(EX833) );
and2 gate( .a(N2235_NOT), .b(EX833), .O(EX834) );
and2 gate( .a(N2228_NOT), .b(p335), .O(EX835) );
and2 gate( .a(N2235), .b(EX835), .O(EX836) );
and2 gate( .a(N2228), .b(p336), .O(EX837) );
and2 gate( .a(N2235), .b(EX837), .O(EX838) );
or2  gate( .a(EX832), .b(EX834), .O(EX839) );
or2  gate( .a(EX836), .b(EX839), .O(EX840) );
or2  gate( .a(EX838), .b(EX840), .O(N2245) );
inv1 gate687( .a(N2236), .O(N2250) );
inv1 gate688( .a(N2240), .O(N2253) );
inv1 gate689( .a(N2244), .O(N2256) );
inv1 gate690( .a(N2237), .O(N2257) );
buf1 gate691( .a(N2237), .O(N2260) );
inv1 gate692( .a(N2241), .O(N2263) );
inv1 gate( .a(N1164),.O(N1164_NOT) );
inv1 gate( .a(N2241),.O(N2241_NOT));
and2 gate( .a(N1164_NOT), .b(p337), .O(EX841) );
and2 gate( .a(N2241_NOT), .b(EX841), .O(EX842) );
and2 gate( .a(N1164), .b(p338), .O(EX843) );
and2 gate( .a(N2241_NOT), .b(EX843), .O(EX844) );
and2 gate( .a(N1164_NOT), .b(p339), .O(EX845) );
and2 gate( .a(N2241), .b(EX845), .O(EX846) );
and2 gate( .a(N1164), .b(p340), .O(EX847) );
and2 gate( .a(N2241), .b(EX847), .O(EX848) );
or2  gate( .a(EX842), .b(EX844), .O(EX849) );
or2  gate( .a(EX846), .b(EX849), .O(EX850) );
or2  gate( .a(EX848), .b(EX850), .O(N2266) );
inv1 gate694( .a(N2245), .O(N2269) );
inv1 gate( .a(N1168),.O(N1168_NOT) );
inv1 gate( .a(N2245),.O(N2245_NOT));
and2 gate( .a(N1168_NOT), .b(p341), .O(EX851) );
and2 gate( .a(N2245_NOT), .b(EX851), .O(EX852) );
and2 gate( .a(N1168), .b(p342), .O(EX853) );
and2 gate( .a(N2245_NOT), .b(EX853), .O(EX854) );
and2 gate( .a(N1168_NOT), .b(p343), .O(EX855) );
and2 gate( .a(N2245), .b(EX855), .O(EX856) );
and2 gate( .a(N1168), .b(p344), .O(EX857) );
and2 gate( .a(N2245), .b(EX857), .O(EX858) );
or2  gate( .a(EX852), .b(EX854), .O(EX859) );
or2  gate( .a(EX856), .b(EX859), .O(EX860) );
or2  gate( .a(EX858), .b(EX860), .O(N2272) );
nand8 gate696( .a(N2067), .b(N2012), .c(N2047), .d(N2250), .e(N899), .f(N2256), .g(N2253), .h(N903), .O(N2279) );
buf1 gate697( .a(N2266), .O(N2286) );
buf1 gate698( .a(N2266), .O(N2297) );
buf1 gate699( .a(N2272), .O(N2315) );
buf1 gate700( .a(N2272), .O(N2326) );
and2 gate701( .a(N2086), .b(N2257), .O(N2340) );
and2 gate702( .a(N2089), .b(N2257), .O(N2353) );
and2 gate703( .a(N2086), .b(N2260), .O(N2361) );
inv1 gate( .a(N2089),.O(N2089_NOT) );
inv1 gate( .a(N2260),.O(N2260_NOT));
and2 gate( .a(N2089_NOT), .b(p345), .O(EX861) );
and2 gate( .a(N2260_NOT), .b(EX861), .O(EX862) );
and2 gate( .a(N2089), .b(p346), .O(EX863) );
and2 gate( .a(N2260_NOT), .b(EX863), .O(EX864) );
and2 gate( .a(N2089_NOT), .b(p347), .O(EX865) );
and2 gate( .a(N2260), .b(EX865), .O(EX866) );
and2 gate( .a(N2089), .b(p348), .O(EX867) );
and2 gate( .a(N2260), .b(EX867), .O(EX868) );
or2  gate( .a(EX862), .b(EX864), .O(EX869) );
or2  gate( .a(EX866), .b(EX869), .O(EX870) );
or2  gate( .a(EX868), .b(EX870), .O(N2375) );
and4 gate705( .a(N338), .b(N2279), .c(N313), .d(N313), .O(N2384) );
and2 gate706( .a(N1163), .b(N2263), .O(N2385) );
inv1 gate( .a(N1164),.O(N1164_NOT) );
inv1 gate( .a(N2263),.O(N2263_NOT));
and2 gate( .a(N1164_NOT), .b(p349), .O(EX871) );
and2 gate( .a(N2263_NOT), .b(EX871), .O(EX872) );
and2 gate( .a(N1164), .b(p350), .O(EX873) );
and2 gate( .a(N2263_NOT), .b(EX873), .O(EX874) );
and2 gate( .a(N1164_NOT), .b(p351), .O(EX875) );
and2 gate( .a(N2263), .b(EX875), .O(EX876) );
and2 gate( .a(N1164), .b(p352), .O(EX877) );
and2 gate( .a(N2263), .b(EX877), .O(EX878) );
or2  gate( .a(EX872), .b(EX874), .O(EX879) );
or2  gate( .a(EX876), .b(EX879), .O(EX880) );
or2  gate( .a(EX878), .b(EX880), .O(N2386) );
and2 gate708( .a(N1167), .b(N2269), .O(N2426) );
and2 gate709( .a(N1168), .b(N2269), .O(N2427) );
nand5 gate710( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2537) );
nand5 gate711( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2540) );
nand5 gate712( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2543) );
nand5 gate713( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2546) );
nand5 gate714( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2549) );
nand5 gate715( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2552) );
nand5 gate716( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2555) );
and5 gate717( .a(N2286), .b(N2315), .c(N2361), .d(N2104), .e(N1171), .O(N2558) );
and5 gate718( .a(N2286), .b(N2315), .c(N2340), .d(N2129), .e(N1171), .O(N2561) );
and5 gate719( .a(N2286), .b(N2315), .c(N2340), .d(N2119), .e(N1171), .O(N2564) );
and5 gate720( .a(N2286), .b(N2315), .c(N2353), .d(N2104), .e(N1171), .O(N2567) );
and5 gate721( .a(N2297), .b(N2315), .c(N2375), .d(N2119), .e(N1188), .O(N2570) );
and5 gate722( .a(N2297), .b(N2326), .c(N2361), .d(N2143), .e(N1188), .O(N2573) );
and5 gate723( .a(N2297), .b(N2326), .c(N2375), .d(N2129), .e(N1188), .O(N2576) );
nand5 gate724( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2594) );
nand5 gate725( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2597) );
nand5 gate726( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2600) );
nand5 gate727( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2603) );
nand5 gate728( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2606) );
nand5 gate729( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2611) );
nand5 gate730( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2614) );
nand5 gate731( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2617) );
nand5 gate732( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2620) );
nand5 gate733( .a(N2297), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2627) );
nand5 gate734( .a(N2386), .b(N2326), .c(N2340), .d(N2104), .e(N926), .O(N2628) );
nand5 gate735( .a(N2386), .b(N2427), .c(N2361), .d(N2104), .e(N926), .O(N2629) );
nand5 gate736( .a(N2386), .b(N2427), .c(N2340), .d(N2129), .e(N926), .O(N2630) );
nand5 gate737( .a(N2386), .b(N2427), .c(N2340), .d(N2119), .e(N926), .O(N2631) );
nand5 gate738( .a(N2386), .b(N2427), .c(N2353), .d(N2104), .e(N926), .O(N2632) );
nand5 gate739( .a(N2386), .b(N2426), .c(N2340), .d(N2104), .e(N926), .O(N2633) );
nand5 gate740( .a(N2385), .b(N2427), .c(N2340), .d(N2104), .e(N926), .O(N2634) );
and5 gate741( .a(N2286), .b(N2427), .c(N2361), .d(N2129), .e(N1171), .O(N2639) );
and5 gate742( .a(N2297), .b(N2427), .c(N2361), .d(N2119), .e(N1171), .O(N2642) );
and5 gate743( .a(N2297), .b(N2427), .c(N2375), .d(N2104), .e(N1171), .O(N2645) );
and5 gate744( .a(N2297), .b(N2427), .c(N2340), .d(N2143), .e(N1171), .O(N2648) );
and5 gate745( .a(N2297), .b(N2427), .c(N2353), .d(N2129), .e(N1188), .O(N2651) );
and5 gate746( .a(N2386), .b(N2326), .c(N2361), .d(N2129), .e(N1188), .O(N2655) );
and5 gate747( .a(N2386), .b(N2326), .c(N2361), .d(N2119), .e(N1188), .O(N2658) );
and5 gate748( .a(N2386), .b(N2326), .c(N2375), .d(N2104), .e(N1188), .O(N2661) );
and5 gate749( .a(N2386), .b(N2326), .c(N2353), .d(N2129), .e(N1188), .O(N2664) );
nand2 gate750( .a(N2558), .b(N534), .O(N2669) );
inv1 gate751( .a(N2558), .O(N2670) );
nand2 gate752( .a(N2561), .b(N535), .O(N2671) );
inv1 gate753( .a(N2561), .O(N2672) );
nand2 gate754( .a(N2564), .b(N536), .O(N2673) );
inv1 gate755( .a(N2564), .O(N2674) );
inv1 gate( .a(N2567),.O(N2567_NOT) );
inv1 gate( .a(N537),.O(N537_NOT));
and2 gate( .a(N2567_NOT), .b(p353), .O(EX881) );
and2 gate( .a(N537_NOT), .b(EX881), .O(EX882) );
and2 gate( .a(N2567), .b(p354), .O(EX883) );
and2 gate( .a(N537_NOT), .b(EX883), .O(EX884) );
and2 gate( .a(N2567_NOT), .b(p355), .O(EX885) );
and2 gate( .a(N537), .b(EX885), .O(EX886) );
and2 gate( .a(N2567), .b(p356), .O(EX887) );
and2 gate( .a(N537), .b(EX887), .O(EX888) );
or2  gate( .a(EX882), .b(EX884), .O(EX889) );
or2  gate( .a(EX886), .b(EX889), .O(EX890) );
or2  gate( .a(EX888), .b(EX890), .O(N2675) );
inv1 gate757( .a(N2567), .O(N2676) );
nand2 gate758( .a(N2570), .b(N543), .O(N2682) );
inv1 gate759( .a(N2570), .O(N2683) );
nand2 gate760( .a(N2573), .b(N548), .O(N2688) );
inv1 gate761( .a(N2573), .O(N2689) );
nand2 gate762( .a(N2576), .b(N549), .O(N2690) );
inv1 gate763( .a(N2576), .O(N2691) );
and8 gate764( .a(N2627), .b(N2628), .c(N2629), .d(N2630), .e(N2631), .f(N2632), .g(N2633), .h(N2634), .O(N2710) );
nand2 gate765( .a(N343), .b(N2670), .O(N2720) );
nand2 gate766( .a(N346), .b(N2672), .O(N2721) );
nand2 gate767( .a(N349), .b(N2674), .O(N2722) );
inv1 gate( .a(N352),.O(N352_NOT) );
inv1 gate( .a(N2676),.O(N2676_NOT));
and2 gate( .a(N352_NOT), .b(p357), .O(EX891) );
and2 gate( .a(N2676_NOT), .b(EX891), .O(EX892) );
and2 gate( .a(N352), .b(p358), .O(EX893) );
and2 gate( .a(N2676_NOT), .b(EX893), .O(EX894) );
and2 gate( .a(N352_NOT), .b(p359), .O(EX895) );
and2 gate( .a(N2676), .b(EX895), .O(EX896) );
and2 gate( .a(N352), .b(p360), .O(EX897) );
and2 gate( .a(N2676), .b(EX897), .O(EX898) );
or2  gate( .a(EX892), .b(EX894), .O(EX899) );
or2  gate( .a(EX896), .b(EX899), .O(EX900) );
or2  gate( .a(EX898), .b(EX900), .O(N2723) );
nand2 gate769( .a(N2639), .b(N538), .O(N2724) );
inv1 gate770( .a(N2639), .O(N2725) );
nand2 gate771( .a(N2642), .b(N539), .O(N2726) );
inv1 gate772( .a(N2642), .O(N2727) );
nand2 gate773( .a(N2645), .b(N540), .O(N2728) );
inv1 gate774( .a(N2645), .O(N2729) );
nand2 gate775( .a(N2648), .b(N541), .O(N2730) );
inv1 gate776( .a(N2648), .O(N2731) );
nand2 gate777( .a(N2651), .b(N542), .O(N2732) );
inv1 gate778( .a(N2651), .O(N2733) );
inv1 gate( .a(N370),.O(N370_NOT) );
inv1 gate( .a(N2683),.O(N2683_NOT));
and2 gate( .a(N370_NOT), .b(p361), .O(EX901) );
and2 gate( .a(N2683_NOT), .b(EX901), .O(EX902) );
and2 gate( .a(N370), .b(p362), .O(EX903) );
and2 gate( .a(N2683_NOT), .b(EX903), .O(EX904) );
and2 gate( .a(N370_NOT), .b(p363), .O(EX905) );
and2 gate( .a(N2683), .b(EX905), .O(EX906) );
and2 gate( .a(N370), .b(p364), .O(EX907) );
and2 gate( .a(N2683), .b(EX907), .O(EX908) );
or2  gate( .a(EX902), .b(EX904), .O(EX909) );
or2  gate( .a(EX906), .b(EX909), .O(EX910) );
or2  gate( .a(EX908), .b(EX910), .O(N2734) );
nand2 gate780( .a(N2655), .b(N544), .O(N2735) );
inv1 gate781( .a(N2655), .O(N2736) );
nand2 gate782( .a(N2658), .b(N545), .O(N2737) );
inv1 gate783( .a(N2658), .O(N2738) );
nand2 gate784( .a(N2661), .b(N546), .O(N2739) );
inv1 gate785( .a(N2661), .O(N2740) );
nand2 gate786( .a(N2664), .b(N547), .O(N2741) );
inv1 gate787( .a(N2664), .O(N2742) );
nand2 gate788( .a(N385), .b(N2689), .O(N2743) );
nand2 gate789( .a(N388), .b(N2691), .O(N2744) );
nand8 gate790( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2745) );
nand8 gate791( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2746) );
and8 gate792( .a(N2537), .b(N2540), .c(N2543), .d(N2546), .e(N2594), .f(N2597), .g(N2600), .h(N2603), .O(N2747) );
and8 gate793( .a(N2606), .b(N2549), .c(N2611), .d(N2614), .e(N2617), .f(N2620), .g(N2552), .h(N2555), .O(N2750) );
nand2 gate794( .a(N2669), .b(N2720), .O(N2753) );
nand2 gate795( .a(N2671), .b(N2721), .O(N2754) );
inv1 gate( .a(N2673),.O(N2673_NOT) );
inv1 gate( .a(N2722),.O(N2722_NOT));
and2 gate( .a(N2673_NOT), .b(p365), .O(EX911) );
and2 gate( .a(N2722_NOT), .b(EX911), .O(EX912) );
and2 gate( .a(N2673), .b(p366), .O(EX913) );
and2 gate( .a(N2722_NOT), .b(EX913), .O(EX914) );
and2 gate( .a(N2673_NOT), .b(p367), .O(EX915) );
and2 gate( .a(N2722), .b(EX915), .O(EX916) );
and2 gate( .a(N2673), .b(p368), .O(EX917) );
and2 gate( .a(N2722), .b(EX917), .O(EX918) );
or2  gate( .a(EX912), .b(EX914), .O(EX919) );
or2  gate( .a(EX916), .b(EX919), .O(EX920) );
or2  gate( .a(EX918), .b(EX920), .O(N2755) );
nand2 gate797( .a(N2675), .b(N2723), .O(N2756) );
nand2 gate798( .a(N355), .b(N2725), .O(N2757) );
nand2 gate799( .a(N358), .b(N2727), .O(N2758) );
inv1 gate( .a(N361),.O(N361_NOT) );
inv1 gate( .a(N2729),.O(N2729_NOT));
and2 gate( .a(N361_NOT), .b(p369), .O(EX921) );
and2 gate( .a(N2729_NOT), .b(EX921), .O(EX922) );
and2 gate( .a(N361), .b(p370), .O(EX923) );
and2 gate( .a(N2729_NOT), .b(EX923), .O(EX924) );
and2 gate( .a(N361_NOT), .b(p371), .O(EX925) );
and2 gate( .a(N2729), .b(EX925), .O(EX926) );
and2 gate( .a(N361), .b(p372), .O(EX927) );
and2 gate( .a(N2729), .b(EX927), .O(EX928) );
or2  gate( .a(EX922), .b(EX924), .O(EX929) );
or2  gate( .a(EX926), .b(EX929), .O(EX930) );
or2  gate( .a(EX928), .b(EX930), .O(N2759) );
inv1 gate( .a(N364),.O(N364_NOT) );
inv1 gate( .a(N2731),.O(N2731_NOT));
and2 gate( .a(N364_NOT), .b(p373), .O(EX931) );
and2 gate( .a(N2731_NOT), .b(EX931), .O(EX932) );
and2 gate( .a(N364), .b(p374), .O(EX933) );
and2 gate( .a(N2731_NOT), .b(EX933), .O(EX934) );
and2 gate( .a(N364_NOT), .b(p375), .O(EX935) );
and2 gate( .a(N2731), .b(EX935), .O(EX936) );
and2 gate( .a(N364), .b(p376), .O(EX937) );
and2 gate( .a(N2731), .b(EX937), .O(EX938) );
or2  gate( .a(EX932), .b(EX934), .O(EX939) );
or2  gate( .a(EX936), .b(EX939), .O(EX940) );
or2  gate( .a(EX938), .b(EX940), .O(N2760) );
nand2 gate802( .a(N367), .b(N2733), .O(N2761) );
nand2 gate803( .a(N2682), .b(N2734), .O(N2762) );
nand2 gate804( .a(N373), .b(N2736), .O(N2763) );
nand2 gate805( .a(N376), .b(N2738), .O(N2764) );
inv1 gate( .a(N379),.O(N379_NOT) );
inv1 gate( .a(N2740),.O(N2740_NOT));
and2 gate( .a(N379_NOT), .b(p377), .O(EX941) );
and2 gate( .a(N2740_NOT), .b(EX941), .O(EX942) );
and2 gate( .a(N379), .b(p378), .O(EX943) );
and2 gate( .a(N2740_NOT), .b(EX943), .O(EX944) );
and2 gate( .a(N379_NOT), .b(p379), .O(EX945) );
and2 gate( .a(N2740), .b(EX945), .O(EX946) );
and2 gate( .a(N379), .b(p380), .O(EX947) );
and2 gate( .a(N2740), .b(EX947), .O(EX948) );
or2  gate( .a(EX942), .b(EX944), .O(EX949) );
or2  gate( .a(EX946), .b(EX949), .O(EX950) );
or2  gate( .a(EX948), .b(EX950), .O(N2765) );
nand2 gate807( .a(N382), .b(N2742), .O(N2766) );
nand2 gate808( .a(N2688), .b(N2743), .O(N2767) );
nand2 gate809( .a(N2690), .b(N2744), .O(N2768) );
and2 gate810( .a(N2745), .b(N275), .O(N2773) );
and2 gate811( .a(N2746), .b(N276), .O(N2776) );
nand2 gate812( .a(N2724), .b(N2757), .O(N2779) );
nand2 gate813( .a(N2726), .b(N2758), .O(N2780) );
nand2 gate814( .a(N2728), .b(N2759), .O(N2781) );
nand2 gate815( .a(N2730), .b(N2760), .O(N2782) );
nand2 gate816( .a(N2732), .b(N2761), .O(N2783) );
nand2 gate817( .a(N2735), .b(N2763), .O(N2784) );
nand2 gate818( .a(N2737), .b(N2764), .O(N2785) );
nand2 gate819( .a(N2739), .b(N2765), .O(N2786) );
nand2 gate820( .a(N2741), .b(N2766), .O(N2787) );
and3 gate821( .a(N2747), .b(N2750), .c(N2710), .O(N2788) );
nand2 gate822( .a(N2747), .b(N2750), .O(N2789) );
and4 gate823( .a(N338), .b(N2279), .c(N99), .d(N2788), .O(N2800) );
nand2 gate824( .a(N2773), .b(N2018), .O(N2807) );
inv1 gate825( .a(N2773), .O(N2808) );
inv1 gate( .a(N2776),.O(N2776_NOT) );
inv1 gate( .a(N2019),.O(N2019_NOT));
and2 gate( .a(N2776_NOT), .b(p381), .O(EX951) );
and2 gate( .a(N2019_NOT), .b(EX951), .O(EX952) );
and2 gate( .a(N2776), .b(p382), .O(EX953) );
and2 gate( .a(N2019_NOT), .b(EX953), .O(EX954) );
and2 gate( .a(N2776_NOT), .b(p383), .O(EX955) );
and2 gate( .a(N2019), .b(EX955), .O(EX956) );
and2 gate( .a(N2776), .b(p384), .O(EX957) );
and2 gate( .a(N2019), .b(EX957), .O(EX958) );
or2  gate( .a(EX952), .b(EX954), .O(EX959) );
or2  gate( .a(EX956), .b(EX959), .O(EX960) );
or2  gate( .a(EX958), .b(EX960), .O(N2809) );
inv1 gate827( .a(N2776), .O(N2810) );
inv1 gate( .a(N2384),.O(N2384_NOT) );
inv1 gate( .a(N2800),.O(N2800_NOT));
and2 gate( .a(N2384_NOT), .b(p385), .O(EX961) );
and2 gate( .a(N2800_NOT), .b(EX961), .O(EX962) );
and2 gate( .a(N2384), .b(p386), .O(EX963) );
and2 gate( .a(N2800_NOT), .b(EX963), .O(EX964) );
and2 gate( .a(N2384_NOT), .b(p387), .O(EX965) );
and2 gate( .a(N2800), .b(EX965), .O(EX966) );
and2 gate( .a(N2384), .b(p388), .O(EX967) );
and2 gate( .a(N2800), .b(EX967), .O(EX968) );
or2  gate( .a(EX962), .b(EX964), .O(EX969) );
or2  gate( .a(EX966), .b(EX969), .O(EX970) );
or2  gate( .a(EX968), .b(EX970), .O(N2811) );
and3 gate829( .a(N897), .b(N283), .c(N2789), .O(N2812) );
and3 gate830( .a(N76), .b(N283), .c(N2789), .O(N2815) );
and3 gate831( .a(N82), .b(N283), .c(N2789), .O(N2818) );
and3 gate832( .a(N85), .b(N283), .c(N2789), .O(N2821) );
and3 gate833( .a(N898), .b(N283), .c(N2789), .O(N2824) );
nand2 gate834( .a(N1965), .b(N2808), .O(N2827) );
nand2 gate835( .a(N1968), .b(N2810), .O(N2828) );
and3 gate836( .a(N79), .b(N283), .c(N2789), .O(N2829) );
nand2 gate837( .a(N2807), .b(N2827), .O(N2843) );
nand2 gate838( .a(N2809), .b(N2828), .O(N2846) );
nand2 gate839( .a(N2812), .b(N2076), .O(N2850) );
nand2 gate840( .a(N2815), .b(N2077), .O(N2851) );
nand2 gate841( .a(N2818), .b(N1915), .O(N2852) );
nand2 gate842( .a(N2821), .b(N1857), .O(N2853) );
nand2 gate843( .a(N2824), .b(N1938), .O(N2854) );
inv1 gate844( .a(N2812), .O(N2857) );
inv1 gate845( .a(N2815), .O(N2858) );
inv1 gate846( .a(N2818), .O(N2859) );
inv1 gate847( .a(N2821), .O(N2860) );
inv1 gate848( .a(N2824), .O(N2861) );
inv1 gate849( .a(N2829), .O(N2862) );
inv1 gate( .a(N2829),.O(N2829_NOT) );
inv1 gate( .a(N1985),.O(N1985_NOT));
and2 gate( .a(N2829_NOT), .b(p389), .O(EX971) );
and2 gate( .a(N1985_NOT), .b(EX971), .O(EX972) );
and2 gate( .a(N2829), .b(p390), .O(EX973) );
and2 gate( .a(N1985_NOT), .b(EX973), .O(EX974) );
and2 gate( .a(N2829_NOT), .b(p391), .O(EX975) );
and2 gate( .a(N1985), .b(EX975), .O(EX976) );
and2 gate( .a(N2829), .b(p392), .O(EX977) );
and2 gate( .a(N1985), .b(EX977), .O(EX978) );
or2  gate( .a(EX972), .b(EX974), .O(EX979) );
or2  gate( .a(EX976), .b(EX979), .O(EX980) );
or2  gate( .a(EX978), .b(EX980), .O(N2863) );
nand2 gate851( .a(N2052), .b(N2857), .O(N2866) );
nand2 gate852( .a(N2055), .b(N2858), .O(N2867) );
inv1 gate( .a(N1866),.O(N1866_NOT) );
inv1 gate( .a(N2859),.O(N2859_NOT));
and2 gate( .a(N1866_NOT), .b(p393), .O(EX981) );
and2 gate( .a(N2859_NOT), .b(EX981), .O(EX982) );
and2 gate( .a(N1866), .b(p394), .O(EX983) );
and2 gate( .a(N2859_NOT), .b(EX983), .O(EX984) );
and2 gate( .a(N1866_NOT), .b(p395), .O(EX985) );
and2 gate( .a(N2859), .b(EX985), .O(EX986) );
and2 gate( .a(N1866), .b(p396), .O(EX987) );
and2 gate( .a(N2859), .b(EX987), .O(EX988) );
or2  gate( .a(EX982), .b(EX984), .O(EX989) );
or2  gate( .a(EX986), .b(EX989), .O(EX990) );
or2  gate( .a(EX988), .b(EX990), .O(N2868) );
nand2 gate854( .a(N1818), .b(N2860), .O(N2869) );
inv1 gate( .a(N1902),.O(N1902_NOT) );
inv1 gate( .a(N2861),.O(N2861_NOT));
and2 gate( .a(N1902_NOT), .b(p397), .O(EX991) );
and2 gate( .a(N2861_NOT), .b(EX991), .O(EX992) );
and2 gate( .a(N1902), .b(p398), .O(EX993) );
and2 gate( .a(N2861_NOT), .b(EX993), .O(EX994) );
and2 gate( .a(N1902_NOT), .b(p399), .O(EX995) );
and2 gate( .a(N2861), .b(EX995), .O(EX996) );
and2 gate( .a(N1902), .b(p400), .O(EX997) );
and2 gate( .a(N2861), .b(EX997), .O(EX998) );
or2  gate( .a(EX992), .b(EX994), .O(EX999) );
or2  gate( .a(EX996), .b(EX999), .O(EX1000) );
or2  gate( .a(EX998), .b(EX1000), .O(N2870) );
inv1 gate( .a(N2843),.O(N2843_NOT) );
inv1 gate( .a(N886),.O(N886_NOT));
and2 gate( .a(N2843_NOT), .b(p401), .O(EX1001) );
and2 gate( .a(N886_NOT), .b(EX1001), .O(EX1002) );
and2 gate( .a(N2843), .b(p402), .O(EX1003) );
and2 gate( .a(N886_NOT), .b(EX1003), .O(EX1004) );
and2 gate( .a(N2843_NOT), .b(p403), .O(EX1005) );
and2 gate( .a(N886), .b(EX1005), .O(EX1006) );
and2 gate( .a(N2843), .b(p404), .O(EX1007) );
and2 gate( .a(N886), .b(EX1007), .O(EX1008) );
or2  gate( .a(EX1002), .b(EX1004), .O(EX1009) );
or2  gate( .a(EX1006), .b(EX1009), .O(EX1010) );
or2  gate( .a(EX1008), .b(EX1010), .O(N2871) );
inv1 gate857( .a(N2843), .O(N2872) );
inv1 gate( .a(N2846),.O(N2846_NOT) );
inv1 gate( .a(N887),.O(N887_NOT));
and2 gate( .a(N2846_NOT), .b(p405), .O(EX1011) );
and2 gate( .a(N887_NOT), .b(EX1011), .O(EX1012) );
and2 gate( .a(N2846), .b(p406), .O(EX1013) );
and2 gate( .a(N887_NOT), .b(EX1013), .O(EX1014) );
and2 gate( .a(N2846_NOT), .b(p407), .O(EX1015) );
and2 gate( .a(N887), .b(EX1015), .O(EX1016) );
and2 gate( .a(N2846), .b(p408), .O(EX1017) );
and2 gate( .a(N887), .b(EX1017), .O(EX1018) );
or2  gate( .a(EX1012), .b(EX1014), .O(EX1019) );
or2  gate( .a(EX1016), .b(EX1019), .O(EX1020) );
or2  gate( .a(EX1018), .b(EX1020), .O(N2873) );
inv1 gate859( .a(N2846), .O(N2874) );
nand2 gate860( .a(N1933), .b(N2862), .O(N2875) );
nand2 gate861( .a(N2866), .b(N2850), .O(N2876) );
nand2 gate862( .a(N2867), .b(N2851), .O(N2877) );
nand2 gate863( .a(N2868), .b(N2852), .O(N2878) );
nand2 gate864( .a(N2869), .b(N2853), .O(N2879) );
nand2 gate865( .a(N2870), .b(N2854), .O(N2880) );
nand2 gate866( .a(N682), .b(N2872), .O(N2881) );
inv1 gate( .a(N685),.O(N685_NOT) );
inv1 gate( .a(N2874),.O(N2874_NOT));
and2 gate( .a(N685_NOT), .b(p409), .O(EX1021) );
and2 gate( .a(N2874_NOT), .b(EX1021), .O(EX1022) );
and2 gate( .a(N685), .b(p410), .O(EX1023) );
and2 gate( .a(N2874_NOT), .b(EX1023), .O(EX1024) );
and2 gate( .a(N685_NOT), .b(p411), .O(EX1025) );
and2 gate( .a(N2874), .b(EX1025), .O(EX1026) );
and2 gate( .a(N685), .b(p412), .O(EX1027) );
and2 gate( .a(N2874), .b(EX1027), .O(EX1028) );
or2  gate( .a(EX1022), .b(EX1024), .O(EX1029) );
or2  gate( .a(EX1026), .b(EX1029), .O(EX1030) );
or2  gate( .a(EX1028), .b(EX1030), .O(N2882) );
nand2 gate868( .a(N2875), .b(N2863), .O(N2883) );
and2 gate869( .a(N2876), .b(N550), .O(N2886) );
and2 gate870( .a(N551), .b(N2877), .O(N2887) );
and2 gate871( .a(N553), .b(N2878), .O(N2888) );
and2 gate872( .a(N2879), .b(N554), .O(N2889) );
and2 gate873( .a(N555), .b(N2880), .O(N2890) );
inv1 gate( .a(N2871),.O(N2871_NOT) );
inv1 gate( .a(N2881),.O(N2881_NOT));
and2 gate( .a(N2871_NOT), .b(p413), .O(EX1031) );
and2 gate( .a(N2881_NOT), .b(EX1031), .O(EX1032) );
and2 gate( .a(N2871), .b(p414), .O(EX1033) );
and2 gate( .a(N2881_NOT), .b(EX1033), .O(EX1034) );
and2 gate( .a(N2871_NOT), .b(p415), .O(EX1035) );
and2 gate( .a(N2881), .b(EX1035), .O(EX1036) );
and2 gate( .a(N2871), .b(p416), .O(EX1037) );
and2 gate( .a(N2881), .b(EX1037), .O(EX1038) );
or2  gate( .a(EX1032), .b(EX1034), .O(EX1039) );
or2  gate( .a(EX1036), .b(EX1039), .O(EX1040) );
or2  gate( .a(EX1038), .b(EX1040), .O(N2891) );
nand2 gate875( .a(N2873), .b(N2882), .O(N2892) );
nand2 gate876( .a(N2883), .b(N1461), .O(N2895) );
inv1 gate877( .a(N2883), .O(N2896) );
nand2 gate878( .a(N1383), .b(N2896), .O(N2897) );
inv1 gate( .a(N2895),.O(N2895_NOT) );
inv1 gate( .a(N2897),.O(N2897_NOT));
and2 gate( .a(N2895_NOT), .b(p417), .O(EX1041) );
and2 gate( .a(N2897_NOT), .b(EX1041), .O(EX1042) );
and2 gate( .a(N2895), .b(p418), .O(EX1043) );
and2 gate( .a(N2897_NOT), .b(EX1043), .O(EX1044) );
and2 gate( .a(N2895_NOT), .b(p419), .O(EX1045) );
and2 gate( .a(N2897), .b(EX1045), .O(EX1046) );
and2 gate( .a(N2895), .b(p420), .O(EX1047) );
and2 gate( .a(N2897), .b(EX1047), .O(EX1048) );
or2  gate( .a(EX1042), .b(EX1044), .O(EX1049) );
or2  gate( .a(EX1046), .b(EX1049), .O(EX1050) );
or2  gate( .a(EX1048), .b(EX1050), .O(N2898) );
and2 gate880( .a(N2898), .b(N552), .O(N2899) );

endmodule
