
module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;

input p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,
        p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,
        p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,
        p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,
        p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,
        p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,
        p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,
        p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,
        p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,
        p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,
        p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,
        p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,
        p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,
        p131,p132,p133,p134,p135,p136,p137,p138,p139,p140,
        p141,p142,p143,p144,p145,p146,p147,p148,p149,p150,
        p151,p152,p153,p154,p155,p156,p157,p158,p159,p160,
        p161,p162,p163,p164,p165,p166,p167,p168,p169,p170,
        p171,p172,p173,p174,p175,p176,p177,p178,p179,p180,
        p181,p182,p183,p184,p185,p186,p187,p188,p189,p190,
        p191,p192,p193,p194,p195,p196,p197,p198,p199,p200,
        p201,p202,p203,p204,p205,p206,p207,p208,p209,p210,
        p211,p212,p213,p214,p215,p216,p217,p218,p219,p220,
        p221,p222,p223,p224,p225,p226,p227,p228,p229,p230,
        p231,p232,p233,p234,p235,p236,p237,p238,p239,p240,
        p241,p242,p243,p244,p245,p246,p247,p248,p249,p250,
        p251,p252,p253,p254,p255,p256;

output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,
     N9_NOT,N13_NOT,N33_NOT,N37_NOT,N65_NOT,N69_NOT,N73_NOT,N77_NOT,N81_NOT,N85_NOT,
     N89_NOT,N93_NOT,N97_NOT,N101_NOT,N113_NOT,N117_NOT,N131_NOT,N137_NOT,N132_NOT,N137_NOT,
     N133_NOT,N137_NOT,N135_NOT,N137_NOT,N5_NOT,N21_NOT,N41_NOT,N57_NOT,N97_NOT,N113_NOT,
     N109_NOT,N125_NOT,N252_NOT,N253_NOT,N256_NOT,N257_NOT,N260_NOT,N261_NOT,N276_NOT,N277_NOT,
     N278_NOT,N279_NOT,N282_NOT,N283_NOT,N286_NOT,N287_NOT,N288_NOT,N289_NOT,N302_NOT,N305_NOT,
     N302_NOT,N308_NOT,N267_NOT,N343_NOT,N268_NOT,N344_NOT,N269_NOT,N345_NOT,N271_NOT,N339_NOT,
     N272_NOT,N340_NOT,N319_NOT,N351_NOT,N321_NOT,N353_NOT,N367_NOT,N620_NOT,N393_NOT,N625_NOT,
     N354_NOT,N630_NOT,N367_NOT,N630_NOT,N380_NOT,N630_NOT,N393_NOT,N630_NOT,N406_NOT,N650_NOT,
     N419_NOT,N650_NOT,N432_NOT,N650_NOT,N445_NOT,N650_NOT,N406_NOT,N655_NOT,N419_NOT,N655_NOT,
     N5_NOT,N693_NOT,N13_NOT,N695_NOT,N17_NOT,N696_NOT,N21_NOT,N697_NOT,N25_NOT,N698_NOT,
     N29_NOT,N699_NOT,N37_NOT,N701_NOT,N41_NOT,N702_NOT,N61_NOT,N707_NOT,N65_NOT,N708_NOT,
     N69_NOT,N709_NOT,N77_NOT,N711_NOT,N89_NOT,N714_NOT,N93_NOT,N715_NOT,N97_NOT,N716_NOT,
     N109_NOT,N719_NOT,N113_NOT,N720_NOT,N117_NOT,N721_NOT,N121_NOT,N722_NOT,EX1,EX2,EX3,EX4,EX5,EX6,EX7,EX8,EX9,EX10,
     EX11,EX12,EX13,EX14,EX15,EX16,EX17,EX18,EX19,EX20,
     EX21,EX22,EX23,EX24,EX25,EX26,EX27,EX28,EX29,EX30,
     EX31,EX32,EX33,EX34,EX35,EX36,EX37,EX38,EX39,EX40,
     EX41,EX42,EX43,EX44,EX45,EX46,EX47,EX48,EX49,EX50,
     EX51,EX52,EX53,EX54,EX55,EX56,EX57,EX58,EX59,EX60,
     EX61,EX62,EX63,EX64,EX65,EX66,EX67,EX68,EX69,EX70,
     EX71,EX72,EX73,EX74,EX75,EX76,EX77,EX78,EX79,EX80,
     EX81,EX82,EX83,EX84,EX85,EX86,EX87,EX88,EX89,EX90,
     EX91,EX92,EX93,EX94,EX95,EX96,EX97,EX98,EX99,EX100,
     EX101,EX102,EX103,EX104,EX105,EX106,EX107,EX108,EX109,EX110,
     EX111,EX112,EX113,EX114,EX115,EX116,EX117,EX118,EX119,EX120,
     EX121,EX122,EX123,EX124,EX125,EX126,EX127,EX128,EX129,EX130,
     EX131,EX132,EX133,EX134,EX135,EX136,EX137,EX138,EX139,EX140,
     EX141,EX142,EX143,EX144,EX145,EX146,EX147,EX148,EX149,EX150,
     EX151,EX152,EX153,EX154,EX155,EX156,EX157,EX158,EX159,EX160,
     EX161,EX162,EX163,EX164,EX165,EX166,EX167,EX168,EX169,EX170,
     EX171,EX172,EX173,EX174,EX175,EX176,EX177,EX178,EX179,EX180,
     EX181,EX182,EX183,EX184,EX185,EX186,EX187,EX188,EX189,EX190,
     EX191,EX192,EX193,EX194,EX195,EX196,EX197,EX198,EX199,EX200,
     EX201,EX202,EX203,EX204,EX205,EX206,EX207,EX208,EX209,EX210,
     EX211,EX212,EX213,EX214,EX215,EX216,EX217,EX218,EX219,EX220,
     EX221,EX222,EX223,EX224,EX225,EX226,EX227,EX228,EX229,EX230,
     EX231,EX232,EX233,EX234,EX235,EX236,EX237,EX238,EX239,EX240,
     EX241,EX242,EX243,EX244,EX245,EX246,EX247,EX248,EX249,EX250,
     EX251,EX252,EX253,EX254,EX255,EX256,EX257,EX258,EX259,EX260,
     EX261,EX262,EX263,EX264,EX265,EX266,EX267,EX268,EX269,EX270,
     EX271,EX272,EX273,EX274,EX275,EX276,EX277,EX278,EX279,EX280,
     EX281,EX282,EX283,EX284,EX285,EX286,EX287,EX288,EX289,EX290,
     EX291,EX292,EX293,EX294,EX295,EX296,EX297,EX298,EX299,EX300,
     EX301,EX302,EX303,EX304,EX305,EX306,EX307,EX308,EX309,EX310,
     EX311,EX312,EX313,EX314,EX315,EX316,EX317,EX318,EX319,EX320,
     EX321,EX322,EX323,EX324,EX325,EX326,EX327,EX328,EX329,EX330,
     EX331,EX332,EX333,EX334,EX335,EX336,EX337,EX338,EX339,EX340,
     EX341,EX342,EX343,EX344,EX345,EX346,EX347,EX348,EX349,EX350,
     EX351,EX352,EX353,EX354,EX355,EX356,EX357,EX358,EX359,EX360,
     EX361,EX362,EX363,EX364,EX365,EX366,EX367,EX368,EX369,EX370,
     EX371,EX372,EX373,EX374,EX375,EX376,EX377,EX378,EX379,EX380,
     EX381,EX382,EX383,EX384,EX385,EX386,EX387,EX388,EX389,EX390,
     EX391,EX392,EX393,EX394,EX395,EX396,EX397,EX398,EX399,EX400,
     EX401,EX402,EX403,EX404,EX405,EX406,EX407,EX408,EX409,EX410,
     EX411,EX412,EX413,EX414,EX415,EX416,EX417,EX418,EX419,EX420,
     EX421,EX422,EX423,EX424,EX425,EX426,EX427,EX428,EX429,EX430,
     EX431,EX432,EX433,EX434,EX435,EX436,EX437,EX438,EX439,EX440,
     EX441,EX442,EX443,EX444,EX445,EX446,EX447,EX448,EX449,EX450,
     EX451,EX452,EX453,EX454,EX455,EX456,EX457,EX458,EX459,EX460,
     EX461,EX462,EX463,EX464,EX465,EX466,EX467,EX468,EX469,EX470,
     EX471,EX472,EX473,EX474,EX475,EX476,EX477,EX478,EX479,EX480,
     EX481,EX482,EX483,EX484,EX485,EX486,EX487,EX488,EX489,EX490,
     EX491,EX492,EX493,EX494,EX495,EX496,EX497,EX498,EX499,EX500,
     EX501,EX502,EX503,EX504,EX505,EX506,EX507,EX508,EX509,EX510,
     EX511,EX512,EX513,EX514,EX515,EX516,EX517,EX518,EX519,EX520,
     EX521,EX522,EX523,EX524,EX525,EX526,EX527,EX528,EX529,EX530,
     EX531,EX532,EX533,EX534,EX535,EX536,EX537,EX538,EX539,EX540,
     EX541,EX542,EX543,EX544,EX545,EX546,EX547,EX548,EX549,EX550,
     EX551,EX552,EX553,EX554,EX555,EX556,EX557,EX558,EX559,EX560,
     EX561,EX562,EX563,EX564,EX565,EX566,EX567,EX568,EX569,EX570,
     EX571,EX572,EX573,EX574,EX575,EX576,EX577,EX578,EX579,EX580,
     EX581,EX582,EX583,EX584,EX585,EX586,EX587,EX588,EX589,EX590,
     EX591,EX592,EX593,EX594,EX595,EX596,EX597,EX598,EX599,EX600,
     EX601,EX602,EX603,EX604,EX605,EX606,EX607,EX608,EX609,EX610,
     EX611,EX612,EX613,EX614,EX615,EX616,EX617,EX618,EX619,EX620,
     EX621,EX622,EX623,EX624,EX625,EX626,EX627,EX628,EX629,EX630,
     EX631,EX632,EX633,EX634,EX635,EX636,EX637,EX638,EX639,EX640;


xor2 gate1( .a(N1), .b(N5), .O(N250) );
inv1 gate( .a(N9),.O(N9_NOT) );
inv1 gate( .a(N13),.O(N13_NOT));
and2 gate( .a(N9_NOT), .b(p1), .O(EX1) );
and2 gate( .a(N13_NOT), .b(EX1), .O(EX2) );
and2 gate( .a(N9), .b(p2), .O(EX3) );
and2 gate( .a(N13_NOT), .b(EX3), .O(EX4) );
and2 gate( .a(N9_NOT), .b(p3), .O(EX5) );
and2 gate( .a(N13), .b(EX5), .O(EX6) );
and2 gate( .a(N9), .b(p4), .O(EX7) );
and2 gate( .a(N13), .b(EX7), .O(EX8) );
or2  gate( .a(EX2), .b(EX4), .O(EX9) );
or2  gate( .a(EX6), .b(EX9), .O(EX10) );
or2  gate( .a(EX8), .b(EX10), .O(N251) );
xor2 gate3( .a(N17), .b(N21), .O(N252) );
xor2 gate4( .a(N25), .b(N29), .O(N253) );
inv1 gate( .a(N33),.O(N33_NOT) );
inv1 gate( .a(N37),.O(N37_NOT));
and2 gate( .a(N33_NOT), .b(p5), .O(EX11) );
and2 gate( .a(N37_NOT), .b(EX11), .O(EX12) );
and2 gate( .a(N33), .b(p6), .O(EX13) );
and2 gate( .a(N37_NOT), .b(EX13), .O(EX14) );
and2 gate( .a(N33_NOT), .b(p7), .O(EX15) );
and2 gate( .a(N37), .b(EX15), .O(EX16) );
and2 gate( .a(N33), .b(p8), .O(EX17) );
and2 gate( .a(N37), .b(EX17), .O(EX18) );
or2  gate( .a(EX12), .b(EX14), .O(EX19) );
or2  gate( .a(EX16), .b(EX19), .O(EX20) );
or2  gate( .a(EX18), .b(EX20), .O(N254) );
xor2 gate6( .a(N41), .b(N45), .O(N255) );
xor2 gate7( .a(N49), .b(N53), .O(N256) );
xor2 gate8( .a(N57), .b(N61), .O(N257) );
inv1 gate( .a(N65),.O(N65_NOT) );
inv1 gate( .a(N69),.O(N69_NOT));
and2 gate( .a(N65_NOT), .b(p9), .O(EX21) );
and2 gate( .a(N69_NOT), .b(EX21), .O(EX22) );
and2 gate( .a(N65), .b(p10), .O(EX23) );
and2 gate( .a(N69_NOT), .b(EX23), .O(EX24) );
and2 gate( .a(N65_NOT), .b(p11), .O(EX25) );
and2 gate( .a(N69), .b(EX25), .O(EX26) );
and2 gate( .a(N65), .b(p12), .O(EX27) );
and2 gate( .a(N69), .b(EX27), .O(EX28) );
or2  gate( .a(EX22), .b(EX24), .O(EX29) );
or2  gate( .a(EX26), .b(EX29), .O(EX30) );
or2  gate( .a(EX28), .b(EX30), .O(N258) );
inv1 gate( .a(N73),.O(N73_NOT) );
inv1 gate( .a(N77),.O(N77_NOT));
and2 gate( .a(N73_NOT), .b(p13), .O(EX31) );
and2 gate( .a(N77_NOT), .b(EX31), .O(EX32) );
and2 gate( .a(N73), .b(p14), .O(EX33) );
and2 gate( .a(N77_NOT), .b(EX33), .O(EX34) );
and2 gate( .a(N73_NOT), .b(p15), .O(EX35) );
and2 gate( .a(N77), .b(EX35), .O(EX36) );
and2 gate( .a(N73), .b(p16), .O(EX37) );
and2 gate( .a(N77), .b(EX37), .O(EX38) );
or2  gate( .a(EX32), .b(EX34), .O(EX39) );
or2  gate( .a(EX36), .b(EX39), .O(EX40) );
or2  gate( .a(EX38), .b(EX40), .O(N259) );
inv1 gate( .a(N81),.O(N81_NOT) );
inv1 gate( .a(N85),.O(N85_NOT));
and2 gate( .a(N81_NOT), .b(p17), .O(EX41) );
and2 gate( .a(N85_NOT), .b(EX41), .O(EX42) );
and2 gate( .a(N81), .b(p18), .O(EX43) );
and2 gate( .a(N85_NOT), .b(EX43), .O(EX44) );
and2 gate( .a(N81_NOT), .b(p19), .O(EX45) );
and2 gate( .a(N85), .b(EX45), .O(EX46) );
and2 gate( .a(N81), .b(p20), .O(EX47) );
and2 gate( .a(N85), .b(EX47), .O(EX48) );
or2  gate( .a(EX42), .b(EX44), .O(EX49) );
or2  gate( .a(EX46), .b(EX49), .O(EX50) );
or2  gate( .a(EX48), .b(EX50), .O(N260) );
inv1 gate( .a(N89),.O(N89_NOT) );
inv1 gate( .a(N93),.O(N93_NOT));
and2 gate( .a(N89_NOT), .b(p21), .O(EX51) );
and2 gate( .a(N93_NOT), .b(EX51), .O(EX52) );
and2 gate( .a(N89), .b(p22), .O(EX53) );
and2 gate( .a(N93_NOT), .b(EX53), .O(EX54) );
and2 gate( .a(N89_NOT), .b(p23), .O(EX55) );
and2 gate( .a(N93), .b(EX55), .O(EX56) );
and2 gate( .a(N89), .b(p24), .O(EX57) );
and2 gate( .a(N93), .b(EX57), .O(EX58) );
or2  gate( .a(EX52), .b(EX54), .O(EX59) );
or2  gate( .a(EX56), .b(EX59), .O(EX60) );
or2  gate( .a(EX58), .b(EX60), .O(N261) );
inv1 gate( .a(N97),.O(N97_NOT) );
inv1 gate( .a(N101),.O(N101_NOT));
and2 gate( .a(N97_NOT), .b(p25), .O(EX61) );
and2 gate( .a(N101_NOT), .b(EX61), .O(EX62) );
and2 gate( .a(N97), .b(p26), .O(EX63) );
and2 gate( .a(N101_NOT), .b(EX63), .O(EX64) );
and2 gate( .a(N97_NOT), .b(p27), .O(EX65) );
and2 gate( .a(N101), .b(EX65), .O(EX66) );
and2 gate( .a(N97), .b(p28), .O(EX67) );
and2 gate( .a(N101), .b(EX67), .O(EX68) );
or2  gate( .a(EX62), .b(EX64), .O(EX69) );
or2  gate( .a(EX66), .b(EX69), .O(EX70) );
or2  gate( .a(EX68), .b(EX70), .O(N262) );
xor2 gate14( .a(N105), .b(N109), .O(N263) );
inv1 gate( .a(N113),.O(N113_NOT) );
inv1 gate( .a(N117),.O(N117_NOT));
and2 gate( .a(N113_NOT), .b(p29), .O(EX71) );
and2 gate( .a(N117_NOT), .b(EX71), .O(EX72) );
and2 gate( .a(N113), .b(p30), .O(EX73) );
and2 gate( .a(N117_NOT), .b(EX73), .O(EX74) );
and2 gate( .a(N113_NOT), .b(p31), .O(EX75) );
and2 gate( .a(N117), .b(EX75), .O(EX76) );
and2 gate( .a(N113), .b(p32), .O(EX77) );
and2 gate( .a(N117), .b(EX77), .O(EX78) );
or2  gate( .a(EX72), .b(EX74), .O(EX79) );
or2  gate( .a(EX76), .b(EX79), .O(EX80) );
or2  gate( .a(EX78), .b(EX80), .O(N264) );
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
inv1 gate( .a(N131),.O(N131_NOT) );
inv1 gate( .a(N137),.O(N137_NOT));
and2 gate( .a(N131_NOT), .b(p33), .O(EX81) );
and2 gate( .a(N137_NOT), .b(EX81), .O(EX82) );
and2 gate( .a(N131), .b(p34), .O(EX83) );
and2 gate( .a(N137_NOT), .b(EX83), .O(EX84) );
and2 gate( .a(N131_NOT), .b(p35), .O(EX85) );
and2 gate( .a(N137), .b(EX85), .O(EX86) );
and2 gate( .a(N131), .b(p36), .O(EX87) );
and2 gate( .a(N137), .b(EX87), .O(EX88) );
or2  gate( .a(EX82), .b(EX84), .O(EX89) );
or2  gate( .a(EX86), .b(EX89), .O(EX90) );
or2  gate( .a(EX88), .b(EX90), .O(N268) );
inv1 gate( .a(N132),.O(N132_NOT) );
inv1 gate( .a(N137),.O(N137_NOT));
and2 gate( .a(N132_NOT), .b(p37), .O(EX91) );
and2 gate( .a(N137_NOT), .b(EX91), .O(EX92) );
and2 gate( .a(N132), .b(p38), .O(EX93) );
and2 gate( .a(N137_NOT), .b(EX93), .O(EX94) );
and2 gate( .a(N132_NOT), .b(p39), .O(EX95) );
and2 gate( .a(N137), .b(EX95), .O(EX96) );
and2 gate( .a(N132), .b(p40), .O(EX97) );
and2 gate( .a(N137), .b(EX97), .O(EX98) );
or2  gate( .a(EX92), .b(EX94), .O(EX99) );
or2  gate( .a(EX96), .b(EX99), .O(EX100) );
or2  gate( .a(EX98), .b(EX100), .O(N269) );
inv1 gate( .a(N133),.O(N133_NOT) );
inv1 gate( .a(N137),.O(N137_NOT));
and2 gate( .a(N133_NOT), .b(p41), .O(EX101) );
and2 gate( .a(N137_NOT), .b(EX101), .O(EX102) );
and2 gate( .a(N133), .b(p42), .O(EX103) );
and2 gate( .a(N137_NOT), .b(EX103), .O(EX104) );
and2 gate( .a(N133_NOT), .b(p43), .O(EX105) );
and2 gate( .a(N137), .b(EX105), .O(EX106) );
and2 gate( .a(N133), .b(p44), .O(EX107) );
and2 gate( .a(N137), .b(EX107), .O(EX108) );
or2  gate( .a(EX102), .b(EX104), .O(EX109) );
or2  gate( .a(EX106), .b(EX109), .O(EX110) );
or2  gate( .a(EX108), .b(EX110), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
inv1 gate( .a(N135),.O(N135_NOT) );
inv1 gate( .a(N137),.O(N137_NOT));
and2 gate( .a(N135_NOT), .b(p45), .O(EX111) );
and2 gate( .a(N137_NOT), .b(EX111), .O(EX112) );
and2 gate( .a(N135), .b(p46), .O(EX113) );
and2 gate( .a(N137_NOT), .b(EX113), .O(EX114) );
and2 gate( .a(N135_NOT), .b(p47), .O(EX115) );
and2 gate( .a(N137), .b(EX115), .O(EX116) );
and2 gate( .a(N135), .b(p48), .O(EX117) );
and2 gate( .a(N137), .b(EX117), .O(EX118) );
or2  gate( .a(EX112), .b(EX114), .O(EX119) );
or2  gate( .a(EX116), .b(EX119), .O(EX120) );
or2  gate( .a(EX118), .b(EX120), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );
xor2 gate26( .a(N33), .b(N49), .O(N275) );
inv1 gate( .a(N5),.O(N5_NOT) );
inv1 gate( .a(N21),.O(N21_NOT));
and2 gate( .a(N5_NOT), .b(p49), .O(EX121) );
and2 gate( .a(N21_NOT), .b(EX121), .O(EX122) );
and2 gate( .a(N5), .b(p50), .O(EX123) );
and2 gate( .a(N21_NOT), .b(EX123), .O(EX124) );
and2 gate( .a(N5_NOT), .b(p51), .O(EX125) );
and2 gate( .a(N21), .b(EX125), .O(EX126) );
and2 gate( .a(N5), .b(p52), .O(EX127) );
and2 gate( .a(N21), .b(EX127), .O(EX128) );
or2  gate( .a(EX122), .b(EX124), .O(EX129) );
or2  gate( .a(EX126), .b(EX129), .O(EX130) );
or2  gate( .a(EX128), .b(EX130), .O(N276) );
xor2 gate28( .a(N37), .b(N53), .O(N277) );
xor2 gate29( .a(N9), .b(N25), .O(N278) );
inv1 gate( .a(N41),.O(N41_NOT) );
inv1 gate( .a(N57),.O(N57_NOT));
and2 gate( .a(N41_NOT), .b(p53), .O(EX131) );
and2 gate( .a(N57_NOT), .b(EX131), .O(EX132) );
and2 gate( .a(N41), .b(p54), .O(EX133) );
and2 gate( .a(N57_NOT), .b(EX133), .O(EX134) );
and2 gate( .a(N41_NOT), .b(p55), .O(EX135) );
and2 gate( .a(N57), .b(EX135), .O(EX136) );
and2 gate( .a(N41), .b(p56), .O(EX137) );
and2 gate( .a(N57), .b(EX137), .O(EX138) );
or2  gate( .a(EX132), .b(EX134), .O(EX139) );
or2  gate( .a(EX136), .b(EX139), .O(EX140) );
or2  gate( .a(EX138), .b(EX140), .O(N279) );
xor2 gate31( .a(N13), .b(N29), .O(N280) );
xor2 gate32( .a(N45), .b(N61), .O(N281) );
xor2 gate33( .a(N65), .b(N81), .O(N282) );
inv1 gate( .a(N97),.O(N97_NOT) );
inv1 gate( .a(N113),.O(N113_NOT));
and2 gate( .a(N97_NOT), .b(p57), .O(EX141) );
and2 gate( .a(N113_NOT), .b(EX141), .O(EX142) );
and2 gate( .a(N97), .b(p58), .O(EX143) );
and2 gate( .a(N113_NOT), .b(EX143), .O(EX144) );
and2 gate( .a(N97_NOT), .b(p59), .O(EX145) );
and2 gate( .a(N113), .b(EX145), .O(EX146) );
and2 gate( .a(N97), .b(p60), .O(EX147) );
and2 gate( .a(N113), .b(EX147), .O(EX148) );
or2  gate( .a(EX142), .b(EX144), .O(EX149) );
or2  gate( .a(EX146), .b(EX149), .O(EX150) );
or2  gate( .a(EX148), .b(EX150), .O(N283) );
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );
xor2 gate37( .a(N73), .b(N89), .O(N286) );
xor2 gate38( .a(N105), .b(N121), .O(N287) );
xor2 gate39( .a(N77), .b(N93), .O(N288) );
inv1 gate( .a(N109),.O(N109_NOT) );
inv1 gate( .a(N125),.O(N125_NOT));
and2 gate( .a(N109_NOT), .b(p61), .O(EX151) );
and2 gate( .a(N125_NOT), .b(EX151), .O(EX152) );
and2 gate( .a(N109), .b(p62), .O(EX153) );
and2 gate( .a(N125_NOT), .b(EX153), .O(EX154) );
and2 gate( .a(N109_NOT), .b(p63), .O(EX155) );
and2 gate( .a(N125), .b(EX155), .O(EX156) );
and2 gate( .a(N109), .b(p64), .O(EX157) );
and2 gate( .a(N125), .b(EX157), .O(EX158) );
or2  gate( .a(EX152), .b(EX154), .O(EX159) );
or2  gate( .a(EX156), .b(EX159), .O(EX160) );
or2  gate( .a(EX158), .b(EX160), .O(N289) );
xor2 gate41( .a(N250), .b(N251), .O(N290) );
inv1 gate( .a(N252),.O(N252_NOT) );
inv1 gate( .a(N253),.O(N253_NOT));
and2 gate( .a(N252_NOT), .b(p65), .O(EX161) );
and2 gate( .a(N253_NOT), .b(EX161), .O(EX162) );
and2 gate( .a(N252), .b(p66), .O(EX163) );
and2 gate( .a(N253_NOT), .b(EX163), .O(EX164) );
and2 gate( .a(N252_NOT), .b(p67), .O(EX165) );
and2 gate( .a(N253), .b(EX165), .O(EX166) );
and2 gate( .a(N252), .b(p68), .O(EX167) );
and2 gate( .a(N253), .b(EX167), .O(EX168) );
or2  gate( .a(EX162), .b(EX164), .O(EX169) );
or2  gate( .a(EX166), .b(EX169), .O(EX170) );
or2  gate( .a(EX168), .b(EX170), .O(N293) );
xor2 gate43( .a(N254), .b(N255), .O(N296) );
inv1 gate( .a(N256),.O(N256_NOT) );
inv1 gate( .a(N257),.O(N257_NOT));
and2 gate( .a(N256_NOT), .b(p69), .O(EX171) );
and2 gate( .a(N257_NOT), .b(EX171), .O(EX172) );
and2 gate( .a(N256), .b(p70), .O(EX173) );
and2 gate( .a(N257_NOT), .b(EX173), .O(EX174) );
and2 gate( .a(N256_NOT), .b(p71), .O(EX175) );
and2 gate( .a(N257), .b(EX175), .O(EX176) );
and2 gate( .a(N256), .b(p72), .O(EX177) );
and2 gate( .a(N257), .b(EX177), .O(EX178) );
or2  gate( .a(EX172), .b(EX174), .O(EX179) );
or2  gate( .a(EX176), .b(EX179), .O(EX180) );
or2  gate( .a(EX178), .b(EX180), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );
inv1 gate( .a(N260),.O(N260_NOT) );
inv1 gate( .a(N261),.O(N261_NOT));
and2 gate( .a(N260_NOT), .b(p73), .O(EX181) );
and2 gate( .a(N261_NOT), .b(EX181), .O(EX182) );
and2 gate( .a(N260), .b(p74), .O(EX183) );
and2 gate( .a(N261_NOT), .b(EX183), .O(EX184) );
and2 gate( .a(N260_NOT), .b(p75), .O(EX185) );
and2 gate( .a(N261), .b(EX185), .O(EX186) );
and2 gate( .a(N260), .b(p76), .O(EX187) );
and2 gate( .a(N261), .b(EX187), .O(EX188) );
or2  gate( .a(EX182), .b(EX184), .O(EX189) );
or2  gate( .a(EX186), .b(EX189), .O(EX190) );
or2  gate( .a(EX188), .b(EX190), .O(N305) );
xor2 gate47( .a(N262), .b(N263), .O(N308) );
xor2 gate48( .a(N264), .b(N265), .O(N311) );
xor2 gate49( .a(N274), .b(N275), .O(N314) );
inv1 gate( .a(N276),.O(N276_NOT) );
inv1 gate( .a(N277),.O(N277_NOT));
and2 gate( .a(N276_NOT), .b(p77), .O(EX191) );
and2 gate( .a(N277_NOT), .b(EX191), .O(EX192) );
and2 gate( .a(N276), .b(p78), .O(EX193) );
and2 gate( .a(N277_NOT), .b(EX193), .O(EX194) );
and2 gate( .a(N276_NOT), .b(p79), .O(EX195) );
and2 gate( .a(N277), .b(EX195), .O(EX196) );
and2 gate( .a(N276), .b(p80), .O(EX197) );
and2 gate( .a(N277), .b(EX197), .O(EX198) );
or2  gate( .a(EX192), .b(EX194), .O(EX199) );
or2  gate( .a(EX196), .b(EX199), .O(EX200) );
or2  gate( .a(EX198), .b(EX200), .O(N315) );
inv1 gate( .a(N278),.O(N278_NOT) );
inv1 gate( .a(N279),.O(N279_NOT));
and2 gate( .a(N278_NOT), .b(p81), .O(EX201) );
and2 gate( .a(N279_NOT), .b(EX201), .O(EX202) );
and2 gate( .a(N278), .b(p82), .O(EX203) );
and2 gate( .a(N279_NOT), .b(EX203), .O(EX204) );
and2 gate( .a(N278_NOT), .b(p83), .O(EX205) );
and2 gate( .a(N279), .b(EX205), .O(EX206) );
and2 gate( .a(N278), .b(p84), .O(EX207) );
and2 gate( .a(N279), .b(EX207), .O(EX208) );
or2  gate( .a(EX202), .b(EX204), .O(EX209) );
or2  gate( .a(EX206), .b(EX209), .O(EX210) );
or2  gate( .a(EX208), .b(EX210), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );
inv1 gate( .a(N282),.O(N282_NOT) );
inv1 gate( .a(N283),.O(N283_NOT));
and2 gate( .a(N282_NOT), .b(p85), .O(EX211) );
and2 gate( .a(N283_NOT), .b(EX211), .O(EX212) );
and2 gate( .a(N282), .b(p86), .O(EX213) );
and2 gate( .a(N283_NOT), .b(EX213), .O(EX214) );
and2 gate( .a(N282_NOT), .b(p87), .O(EX215) );
and2 gate( .a(N283), .b(EX215), .O(EX216) );
and2 gate( .a(N282), .b(p88), .O(EX217) );
and2 gate( .a(N283), .b(EX217), .O(EX218) );
or2  gate( .a(EX212), .b(EX214), .O(EX219) );
or2  gate( .a(EX216), .b(EX219), .O(EX220) );
or2  gate( .a(EX218), .b(EX220), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );
inv1 gate( .a(N286),.O(N286_NOT) );
inv1 gate( .a(N287),.O(N287_NOT));
and2 gate( .a(N286_NOT), .b(p89), .O(EX221) );
and2 gate( .a(N287_NOT), .b(EX221), .O(EX222) );
and2 gate( .a(N286), .b(p90), .O(EX223) );
and2 gate( .a(N287_NOT), .b(EX223), .O(EX224) );
and2 gate( .a(N286_NOT), .b(p91), .O(EX225) );
and2 gate( .a(N287), .b(EX225), .O(EX226) );
and2 gate( .a(N286), .b(p92), .O(EX227) );
and2 gate( .a(N287), .b(EX227), .O(EX228) );
or2  gate( .a(EX222), .b(EX224), .O(EX229) );
or2  gate( .a(EX226), .b(EX229), .O(EX230) );
or2  gate( .a(EX228), .b(EX230), .O(N320) );
inv1 gate( .a(N288),.O(N288_NOT) );
inv1 gate( .a(N289),.O(N289_NOT));
and2 gate( .a(N288_NOT), .b(p93), .O(EX231) );
and2 gate( .a(N289_NOT), .b(EX231), .O(EX232) );
and2 gate( .a(N288), .b(p94), .O(EX233) );
and2 gate( .a(N289_NOT), .b(EX233), .O(EX234) );
and2 gate( .a(N288_NOT), .b(p95), .O(EX235) );
and2 gate( .a(N289), .b(EX235), .O(EX236) );
and2 gate( .a(N288), .b(p96), .O(EX237) );
and2 gate( .a(N289), .b(EX237), .O(EX238) );
or2  gate( .a(EX232), .b(EX234), .O(EX239) );
or2  gate( .a(EX236), .b(EX239), .O(EX240) );
or2  gate( .a(EX238), .b(EX240), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );
xor2 gate58( .a(N296), .b(N299), .O(N339) );
xor2 gate59( .a(N290), .b(N296), .O(N340) );
xor2 gate60( .a(N293), .b(N299), .O(N341) );
inv1 gate( .a(N302),.O(N302_NOT) );
inv1 gate( .a(N305),.O(N305_NOT));
and2 gate( .a(N302_NOT), .b(p97), .O(EX241) );
and2 gate( .a(N305_NOT), .b(EX241), .O(EX242) );
and2 gate( .a(N302), .b(p98), .O(EX243) );
and2 gate( .a(N305_NOT), .b(EX243), .O(EX244) );
and2 gate( .a(N302_NOT), .b(p99), .O(EX245) );
and2 gate( .a(N305), .b(EX245), .O(EX246) );
and2 gate( .a(N302), .b(p100), .O(EX247) );
and2 gate( .a(N305), .b(EX247), .O(EX248) );
or2  gate( .a(EX242), .b(EX244), .O(EX249) );
or2  gate( .a(EX246), .b(EX249), .O(EX250) );
or2  gate( .a(EX248), .b(EX250), .O(N342) );
xor2 gate62( .a(N308), .b(N311), .O(N343) );
inv1 gate( .a(N302),.O(N302_NOT) );
inv1 gate( .a(N308),.O(N308_NOT));
and2 gate( .a(N302_NOT), .b(p101), .O(EX251) );
and2 gate( .a(N308_NOT), .b(EX251), .O(EX252) );
and2 gate( .a(N302), .b(p102), .O(EX253) );
and2 gate( .a(N308_NOT), .b(EX253), .O(EX254) );
and2 gate( .a(N302_NOT), .b(p103), .O(EX255) );
and2 gate( .a(N308), .b(EX255), .O(EX256) );
and2 gate( .a(N302), .b(p104), .O(EX257) );
and2 gate( .a(N308), .b(EX257), .O(EX258) );
or2  gate( .a(EX252), .b(EX254), .O(EX259) );
or2  gate( .a(EX256), .b(EX259), .O(EX260) );
or2  gate( .a(EX258), .b(EX260), .O(N344) );
xor2 gate64( .a(N305), .b(N311), .O(N345) );
xor2 gate65( .a(N266), .b(N342), .O(N346) );
inv1 gate( .a(N267),.O(N267_NOT) );
inv1 gate( .a(N343),.O(N343_NOT));
and2 gate( .a(N267_NOT), .b(p105), .O(EX261) );
and2 gate( .a(N343_NOT), .b(EX261), .O(EX262) );
and2 gate( .a(N267), .b(p106), .O(EX263) );
and2 gate( .a(N343_NOT), .b(EX263), .O(EX264) );
and2 gate( .a(N267_NOT), .b(p107), .O(EX265) );
and2 gate( .a(N343), .b(EX265), .O(EX266) );
and2 gate( .a(N267), .b(p108), .O(EX267) );
and2 gate( .a(N343), .b(EX267), .O(EX268) );
or2  gate( .a(EX262), .b(EX264), .O(EX269) );
or2  gate( .a(EX266), .b(EX269), .O(EX270) );
or2  gate( .a(EX268), .b(EX270), .O(N347) );
inv1 gate( .a(N268),.O(N268_NOT) );
inv1 gate( .a(N344),.O(N344_NOT));
and2 gate( .a(N268_NOT), .b(p109), .O(EX271) );
and2 gate( .a(N344_NOT), .b(EX271), .O(EX272) );
and2 gate( .a(N268), .b(p110), .O(EX273) );
and2 gate( .a(N344_NOT), .b(EX273), .O(EX274) );
and2 gate( .a(N268_NOT), .b(p111), .O(EX275) );
and2 gate( .a(N344), .b(EX275), .O(EX276) );
and2 gate( .a(N268), .b(p112), .O(EX277) );
and2 gate( .a(N344), .b(EX277), .O(EX278) );
or2  gate( .a(EX272), .b(EX274), .O(EX279) );
or2  gate( .a(EX276), .b(EX279), .O(EX280) );
or2  gate( .a(EX278), .b(EX280), .O(N348) );
inv1 gate( .a(N269),.O(N269_NOT) );
inv1 gate( .a(N345),.O(N345_NOT));
and2 gate( .a(N269_NOT), .b(p113), .O(EX281) );
and2 gate( .a(N345_NOT), .b(EX281), .O(EX282) );
and2 gate( .a(N269), .b(p114), .O(EX283) );
and2 gate( .a(N345_NOT), .b(EX283), .O(EX284) );
and2 gate( .a(N269_NOT), .b(p115), .O(EX285) );
and2 gate( .a(N345), .b(EX285), .O(EX286) );
and2 gate( .a(N269), .b(p116), .O(EX287) );
and2 gate( .a(N345), .b(EX287), .O(EX288) );
or2  gate( .a(EX282), .b(EX284), .O(EX289) );
or2  gate( .a(EX286), .b(EX289), .O(EX290) );
or2  gate( .a(EX288), .b(EX290), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );
inv1 gate( .a(N271),.O(N271_NOT) );
inv1 gate( .a(N339),.O(N339_NOT));
and2 gate( .a(N271_NOT), .b(p117), .O(EX291) );
and2 gate( .a(N339_NOT), .b(EX291), .O(EX292) );
and2 gate( .a(N271), .b(p118), .O(EX293) );
and2 gate( .a(N339_NOT), .b(EX293), .O(EX294) );
and2 gate( .a(N271_NOT), .b(p119), .O(EX295) );
and2 gate( .a(N339), .b(EX295), .O(EX296) );
and2 gate( .a(N271), .b(p120), .O(EX297) );
and2 gate( .a(N339), .b(EX297), .O(EX298) );
or2  gate( .a(EX292), .b(EX294), .O(EX299) );
or2  gate( .a(EX296), .b(EX299), .O(EX300) );
or2  gate( .a(EX298), .b(EX300), .O(N351) );
inv1 gate( .a(N272),.O(N272_NOT) );
inv1 gate( .a(N340),.O(N340_NOT));
and2 gate( .a(N272_NOT), .b(p121), .O(EX301) );
and2 gate( .a(N340_NOT), .b(EX301), .O(EX302) );
and2 gate( .a(N272), .b(p122), .O(EX303) );
and2 gate( .a(N340_NOT), .b(EX303), .O(EX304) );
and2 gate( .a(N272_NOT), .b(p123), .O(EX305) );
and2 gate( .a(N340), .b(EX305), .O(EX306) );
and2 gate( .a(N272), .b(p124), .O(EX307) );
and2 gate( .a(N340), .b(EX307), .O(EX308) );
or2  gate( .a(EX302), .b(EX304), .O(EX309) );
or2  gate( .a(EX306), .b(EX309), .O(EX310) );
or2  gate( .a(EX308), .b(EX310), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );
xor2 gate74( .a(N315), .b(N347), .O(N367) );
xor2 gate75( .a(N316), .b(N348), .O(N380) );
xor2 gate76( .a(N317), .b(N349), .O(N393) );
xor2 gate77( .a(N318), .b(N350), .O(N406) );
inv1 gate( .a(N319),.O(N319_NOT) );
inv1 gate( .a(N351),.O(N351_NOT));
and2 gate( .a(N319_NOT), .b(p125), .O(EX311) );
and2 gate( .a(N351_NOT), .b(EX311), .O(EX312) );
and2 gate( .a(N319), .b(p126), .O(EX313) );
and2 gate( .a(N351_NOT), .b(EX313), .O(EX314) );
and2 gate( .a(N319_NOT), .b(p127), .O(EX315) );
and2 gate( .a(N351), .b(EX315), .O(EX316) );
and2 gate( .a(N319), .b(p128), .O(EX317) );
and2 gate( .a(N351), .b(EX317), .O(EX318) );
or2  gate( .a(EX312), .b(EX314), .O(EX319) );
or2  gate( .a(EX316), .b(EX319), .O(EX320) );
or2  gate( .a(EX318), .b(EX320), .O(N419) );
xor2 gate79( .a(N320), .b(N352), .O(N432) );
inv1 gate( .a(N321),.O(N321_NOT) );
inv1 gate( .a(N353),.O(N353_NOT));
and2 gate( .a(N321_NOT), .b(p129), .O(EX321) );
and2 gate( .a(N353_NOT), .b(EX321), .O(EX322) );
and2 gate( .a(N321), .b(p130), .O(EX323) );
and2 gate( .a(N353_NOT), .b(EX323), .O(EX324) );
and2 gate( .a(N321_NOT), .b(p131), .O(EX325) );
and2 gate( .a(N353), .b(EX325), .O(EX326) );
and2 gate( .a(N321), .b(p132), .O(EX327) );
and2 gate( .a(N353), .b(EX327), .O(EX328) );
or2  gate( .a(EX322), .b(EX324), .O(EX329) );
or2  gate( .a(EX326), .b(EX329), .O(EX330) );
or2  gate( .a(EX328), .b(EX330), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
inv1 gate( .a(N367),.O(N367_NOT) );
inv1 gate( .a(N620),.O(N620_NOT));
and2 gate( .a(N367_NOT), .b(p133), .O(EX331) );
and2 gate( .a(N620_NOT), .b(EX331), .O(EX332) );
and2 gate( .a(N367), .b(p134), .O(EX333) );
and2 gate( .a(N620_NOT), .b(EX333), .O(EX334) );
and2 gate( .a(N367_NOT), .b(p135), .O(EX335) );
and2 gate( .a(N620), .b(EX335), .O(EX336) );
and2 gate( .a(N367), .b(p136), .O(EX337) );
and2 gate( .a(N620), .b(EX337), .O(EX338) );
or2  gate( .a(EX332), .b(EX334), .O(EX339) );
or2  gate( .a(EX336), .b(EX339), .O(EX340) );
or2  gate( .a(EX338), .b(EX340), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
inv1 gate( .a(N393),.O(N393_NOT) );
inv1 gate( .a(N625),.O(N625_NOT));
and2 gate( .a(N393_NOT), .b(p137), .O(EX341) );
and2 gate( .a(N625_NOT), .b(EX341), .O(EX342) );
and2 gate( .a(N393), .b(p138), .O(EX343) );
and2 gate( .a(N625_NOT), .b(EX343), .O(EX344) );
and2 gate( .a(N393_NOT), .b(p139), .O(EX345) );
and2 gate( .a(N625), .b(EX345), .O(EX346) );
and2 gate( .a(N393), .b(p140), .O(EX347) );
and2 gate( .a(N625), .b(EX347), .O(EX348) );
or2  gate( .a(EX342), .b(EX344), .O(EX349) );
or2  gate( .a(EX346), .b(EX349), .O(EX350) );
or2  gate( .a(EX348), .b(EX350), .O(N699) );
inv1 gate( .a(N354),.O(N354_NOT) );
inv1 gate( .a(N630),.O(N630_NOT));
and2 gate( .a(N354_NOT), .b(p141), .O(EX351) );
and2 gate( .a(N630_NOT), .b(EX351), .O(EX352) );
and2 gate( .a(N354), .b(p142), .O(EX353) );
and2 gate( .a(N630_NOT), .b(EX353), .O(EX354) );
and2 gate( .a(N354_NOT), .b(p143), .O(EX355) );
and2 gate( .a(N630), .b(EX355), .O(EX356) );
and2 gate( .a(N354), .b(p144), .O(EX357) );
and2 gate( .a(N630), .b(EX357), .O(EX358) );
or2  gate( .a(EX352), .b(EX354), .O(EX359) );
or2  gate( .a(EX356), .b(EX359), .O(EX360) );
or2  gate( .a(EX358), .b(EX360), .O(N700) );
inv1 gate( .a(N367),.O(N367_NOT) );
inv1 gate( .a(N630),.O(N630_NOT));
and2 gate( .a(N367_NOT), .b(p145), .O(EX361) );
and2 gate( .a(N630_NOT), .b(EX361), .O(EX362) );
and2 gate( .a(N367), .b(p146), .O(EX363) );
and2 gate( .a(N630_NOT), .b(EX363), .O(EX364) );
and2 gate( .a(N367_NOT), .b(p147), .O(EX365) );
and2 gate( .a(N630), .b(EX365), .O(EX366) );
and2 gate( .a(N367), .b(p148), .O(EX367) );
and2 gate( .a(N630), .b(EX367), .O(EX368) );
or2  gate( .a(EX362), .b(EX364), .O(EX369) );
or2  gate( .a(EX366), .b(EX369), .O(EX370) );
or2  gate( .a(EX368), .b(EX370), .O(N701) );
inv1 gate( .a(N380),.O(N380_NOT) );
inv1 gate( .a(N630),.O(N630_NOT));
and2 gate( .a(N380_NOT), .b(p149), .O(EX371) );
and2 gate( .a(N630_NOT), .b(EX371), .O(EX372) );
and2 gate( .a(N380), .b(p150), .O(EX373) );
and2 gate( .a(N630_NOT), .b(EX373), .O(EX374) );
and2 gate( .a(N380_NOT), .b(p151), .O(EX375) );
and2 gate( .a(N630), .b(EX375), .O(EX376) );
and2 gate( .a(N380), .b(p152), .O(EX377) );
and2 gate( .a(N630), .b(EX377), .O(EX378) );
or2  gate( .a(EX372), .b(EX374), .O(EX379) );
or2  gate( .a(EX376), .b(EX379), .O(EX380) );
or2  gate( .a(EX378), .b(EX380), .O(N702) );
inv1 gate( .a(N393),.O(N393_NOT) );
inv1 gate( .a(N630),.O(N630_NOT));
and2 gate( .a(N393_NOT), .b(p153), .O(EX381) );
and2 gate( .a(N630_NOT), .b(EX381), .O(EX382) );
and2 gate( .a(N393), .b(p154), .O(EX383) );
and2 gate( .a(N630_NOT), .b(EX383), .O(EX384) );
and2 gate( .a(N393_NOT), .b(p155), .O(EX385) );
and2 gate( .a(N630), .b(EX385), .O(EX386) );
and2 gate( .a(N393), .b(p156), .O(EX387) );
and2 gate( .a(N630), .b(EX387), .O(EX388) );
or2  gate( .a(EX382), .b(EX384), .O(EX389) );
or2  gate( .a(EX386), .b(EX389), .O(EX390) );
or2  gate( .a(EX388), .b(EX390), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
inv1 gate( .a(N406),.O(N406_NOT) );
inv1 gate( .a(N650),.O(N650_NOT));
and2 gate( .a(N406_NOT), .b(p157), .O(EX391) );
and2 gate( .a(N650_NOT), .b(EX391), .O(EX392) );
and2 gate( .a(N406), .b(p158), .O(EX393) );
and2 gate( .a(N650_NOT), .b(EX393), .O(EX394) );
and2 gate( .a(N406_NOT), .b(p159), .O(EX395) );
and2 gate( .a(N650), .b(EX395), .O(EX396) );
and2 gate( .a(N406), .b(p160), .O(EX397) );
and2 gate( .a(N650), .b(EX397), .O(EX398) );
or2  gate( .a(EX392), .b(EX394), .O(EX399) );
or2  gate( .a(EX396), .b(EX399), .O(EX400) );
or2  gate( .a(EX398), .b(EX400), .O(N716) );
inv1 gate( .a(N419),.O(N419_NOT) );
inv1 gate( .a(N650),.O(N650_NOT));
and2 gate( .a(N419_NOT), .b(p161), .O(EX401) );
and2 gate( .a(N650_NOT), .b(EX401), .O(EX402) );
and2 gate( .a(N419), .b(p162), .O(EX403) );
and2 gate( .a(N650_NOT), .b(EX403), .O(EX404) );
and2 gate( .a(N419_NOT), .b(p163), .O(EX405) );
and2 gate( .a(N650), .b(EX405), .O(EX406) );
and2 gate( .a(N419), .b(p164), .O(EX407) );
and2 gate( .a(N650), .b(EX407), .O(EX408) );
or2  gate( .a(EX402), .b(EX404), .O(EX409) );
or2  gate( .a(EX406), .b(EX409), .O(EX410) );
or2  gate( .a(EX408), .b(EX410), .O(N717) );
inv1 gate( .a(N432),.O(N432_NOT) );
inv1 gate( .a(N650),.O(N650_NOT));
and2 gate( .a(N432_NOT), .b(p165), .O(EX411) );
and2 gate( .a(N650_NOT), .b(EX411), .O(EX412) );
and2 gate( .a(N432), .b(p166), .O(EX413) );
and2 gate( .a(N650_NOT), .b(EX413), .O(EX414) );
and2 gate( .a(N432_NOT), .b(p167), .O(EX415) );
and2 gate( .a(N650), .b(EX415), .O(EX416) );
and2 gate( .a(N432), .b(p168), .O(EX417) );
and2 gate( .a(N650), .b(EX417), .O(EX418) );
or2  gate( .a(EX412), .b(EX414), .O(EX419) );
or2  gate( .a(EX416), .b(EX419), .O(EX420) );
or2  gate( .a(EX418), .b(EX420), .O(N718) );
inv1 gate( .a(N445),.O(N445_NOT) );
inv1 gate( .a(N650),.O(N650_NOT));
and2 gate( .a(N445_NOT), .b(p169), .O(EX421) );
and2 gate( .a(N650_NOT), .b(EX421), .O(EX422) );
and2 gate( .a(N445), .b(p170), .O(EX423) );
and2 gate( .a(N650_NOT), .b(EX423), .O(EX424) );
and2 gate( .a(N445_NOT), .b(p171), .O(EX425) );
and2 gate( .a(N650), .b(EX425), .O(EX426) );
and2 gate( .a(N445), .b(p172), .O(EX427) );
and2 gate( .a(N650), .b(EX427), .O(EX428) );
or2  gate( .a(EX422), .b(EX424), .O(EX429) );
or2  gate( .a(EX426), .b(EX429), .O(EX430) );
or2  gate( .a(EX428), .b(EX430), .O(N719) );
inv1 gate( .a(N406),.O(N406_NOT) );
inv1 gate( .a(N655),.O(N655_NOT));
and2 gate( .a(N406_NOT), .b(p173), .O(EX431) );
and2 gate( .a(N655_NOT), .b(EX431), .O(EX432) );
and2 gate( .a(N406), .b(p174), .O(EX433) );
and2 gate( .a(N655_NOT), .b(EX433), .O(EX434) );
and2 gate( .a(N406_NOT), .b(p175), .O(EX435) );
and2 gate( .a(N655), .b(EX435), .O(EX436) );
and2 gate( .a(N406), .b(p176), .O(EX437) );
and2 gate( .a(N655), .b(EX437), .O(EX438) );
or2  gate( .a(EX432), .b(EX434), .O(EX439) );
or2  gate( .a(EX436), .b(EX439), .O(EX440) );
or2  gate( .a(EX438), .b(EX440), .O(N720) );
inv1 gate( .a(N419),.O(N419_NOT) );
inv1 gate( .a(N655),.O(N655_NOT));
and2 gate( .a(N419_NOT), .b(p177), .O(EX441) );
and2 gate( .a(N655_NOT), .b(EX441), .O(EX442) );
and2 gate( .a(N419), .b(p178), .O(EX443) );
and2 gate( .a(N655_NOT), .b(EX443), .O(EX444) );
and2 gate( .a(N419_NOT), .b(p179), .O(EX445) );
and2 gate( .a(N655), .b(EX445), .O(EX446) );
and2 gate( .a(N419), .b(p180), .O(EX447) );
and2 gate( .a(N655), .b(EX447), .O(EX448) );
or2  gate( .a(EX442), .b(EX444), .O(EX449) );
or2  gate( .a(EX446), .b(EX449), .O(EX450) );
or2  gate( .a(EX448), .b(EX450), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );
inv1 gate( .a(N5),.O(N5_NOT) );
inv1 gate( .a(N693),.O(N693_NOT));
and2 gate( .a(N5_NOT), .b(p181), .O(EX451) );
and2 gate( .a(N693_NOT), .b(EX451), .O(EX452) );
and2 gate( .a(N5), .b(p182), .O(EX453) );
and2 gate( .a(N693_NOT), .b(EX453), .O(EX454) );
and2 gate( .a(N5_NOT), .b(p183), .O(EX455) );
and2 gate( .a(N693), .b(EX455), .O(EX456) );
and2 gate( .a(N5), .b(p184), .O(EX457) );
and2 gate( .a(N693), .b(EX457), .O(EX458) );
or2  gate( .a(EX452), .b(EX454), .O(EX459) );
or2  gate( .a(EX456), .b(EX459), .O(EX460) );
or2  gate( .a(EX458), .b(EX460), .O(N725) );
xor2 gate173( .a(N9), .b(N694), .O(N726) );
inv1 gate( .a(N13),.O(N13_NOT) );
inv1 gate( .a(N695),.O(N695_NOT));
and2 gate( .a(N13_NOT), .b(p185), .O(EX461) );
and2 gate( .a(N695_NOT), .b(EX461), .O(EX462) );
and2 gate( .a(N13), .b(p186), .O(EX463) );
and2 gate( .a(N695_NOT), .b(EX463), .O(EX464) );
and2 gate( .a(N13_NOT), .b(p187), .O(EX465) );
and2 gate( .a(N695), .b(EX465), .O(EX466) );
and2 gate( .a(N13), .b(p188), .O(EX467) );
and2 gate( .a(N695), .b(EX467), .O(EX468) );
or2  gate( .a(EX462), .b(EX464), .O(EX469) );
or2  gate( .a(EX466), .b(EX469), .O(EX470) );
or2  gate( .a(EX468), .b(EX470), .O(N727) );
inv1 gate( .a(N17),.O(N17_NOT) );
inv1 gate( .a(N696),.O(N696_NOT));
and2 gate( .a(N17_NOT), .b(p189), .O(EX471) );
and2 gate( .a(N696_NOT), .b(EX471), .O(EX472) );
and2 gate( .a(N17), .b(p190), .O(EX473) );
and2 gate( .a(N696_NOT), .b(EX473), .O(EX474) );
and2 gate( .a(N17_NOT), .b(p191), .O(EX475) );
and2 gate( .a(N696), .b(EX475), .O(EX476) );
and2 gate( .a(N17), .b(p192), .O(EX477) );
and2 gate( .a(N696), .b(EX477), .O(EX478) );
or2  gate( .a(EX472), .b(EX474), .O(EX479) );
or2  gate( .a(EX476), .b(EX479), .O(EX480) );
or2  gate( .a(EX478), .b(EX480), .O(N728) );
inv1 gate( .a(N21),.O(N21_NOT) );
inv1 gate( .a(N697),.O(N697_NOT));
and2 gate( .a(N21_NOT), .b(p193), .O(EX481) );
and2 gate( .a(N697_NOT), .b(EX481), .O(EX482) );
and2 gate( .a(N21), .b(p194), .O(EX483) );
and2 gate( .a(N697_NOT), .b(EX483), .O(EX484) );
and2 gate( .a(N21_NOT), .b(p195), .O(EX485) );
and2 gate( .a(N697), .b(EX485), .O(EX486) );
and2 gate( .a(N21), .b(p196), .O(EX487) );
and2 gate( .a(N697), .b(EX487), .O(EX488) );
or2  gate( .a(EX482), .b(EX484), .O(EX489) );
or2  gate( .a(EX486), .b(EX489), .O(EX490) );
or2  gate( .a(EX488), .b(EX490), .O(N729) );
inv1 gate( .a(N25),.O(N25_NOT) );
inv1 gate( .a(N698),.O(N698_NOT));
and2 gate( .a(N25_NOT), .b(p197), .O(EX491) );
and2 gate( .a(N698_NOT), .b(EX491), .O(EX492) );
and2 gate( .a(N25), .b(p198), .O(EX493) );
and2 gate( .a(N698_NOT), .b(EX493), .O(EX494) );
and2 gate( .a(N25_NOT), .b(p199), .O(EX495) );
and2 gate( .a(N698), .b(EX495), .O(EX496) );
and2 gate( .a(N25), .b(p200), .O(EX497) );
and2 gate( .a(N698), .b(EX497), .O(EX498) );
or2  gate( .a(EX492), .b(EX494), .O(EX499) );
or2  gate( .a(EX496), .b(EX499), .O(EX500) );
or2  gate( .a(EX498), .b(EX500), .O(N730) );
inv1 gate( .a(N29),.O(N29_NOT) );
inv1 gate( .a(N699),.O(N699_NOT));
and2 gate( .a(N29_NOT), .b(p201), .O(EX501) );
and2 gate( .a(N699_NOT), .b(EX501), .O(EX502) );
and2 gate( .a(N29), .b(p202), .O(EX503) );
and2 gate( .a(N699_NOT), .b(EX503), .O(EX504) );
and2 gate( .a(N29_NOT), .b(p203), .O(EX505) );
and2 gate( .a(N699), .b(EX505), .O(EX506) );
and2 gate( .a(N29), .b(p204), .O(EX507) );
and2 gate( .a(N699), .b(EX507), .O(EX508) );
or2  gate( .a(EX502), .b(EX504), .O(EX509) );
or2  gate( .a(EX506), .b(EX509), .O(EX510) );
or2  gate( .a(EX508), .b(EX510), .O(N731) );
xor2 gate179( .a(N33), .b(N700), .O(N732) );
inv1 gate( .a(N37),.O(N37_NOT) );
inv1 gate( .a(N701),.O(N701_NOT));
and2 gate( .a(N37_NOT), .b(p205), .O(EX511) );
and2 gate( .a(N701_NOT), .b(EX511), .O(EX512) );
and2 gate( .a(N37), .b(p206), .O(EX513) );
and2 gate( .a(N701_NOT), .b(EX513), .O(EX514) );
and2 gate( .a(N37_NOT), .b(p207), .O(EX515) );
and2 gate( .a(N701), .b(EX515), .O(EX516) );
and2 gate( .a(N37), .b(p208), .O(EX517) );
and2 gate( .a(N701), .b(EX517), .O(EX518) );
or2  gate( .a(EX512), .b(EX514), .O(EX519) );
or2  gate( .a(EX516), .b(EX519), .O(EX520) );
or2  gate( .a(EX518), .b(EX520), .O(N733) );
inv1 gate( .a(N41),.O(N41_NOT) );
inv1 gate( .a(N702),.O(N702_NOT));
and2 gate( .a(N41_NOT), .b(p209), .O(EX521) );
and2 gate( .a(N702_NOT), .b(EX521), .O(EX522) );
and2 gate( .a(N41), .b(p210), .O(EX523) );
and2 gate( .a(N702_NOT), .b(EX523), .O(EX524) );
and2 gate( .a(N41_NOT), .b(p211), .O(EX525) );
and2 gate( .a(N702), .b(EX525), .O(EX526) );
and2 gate( .a(N41), .b(p212), .O(EX527) );
and2 gate( .a(N702), .b(EX527), .O(EX528) );
or2  gate( .a(EX522), .b(EX524), .O(EX529) );
or2  gate( .a(EX526), .b(EX529), .O(EX530) );
or2  gate( .a(EX528), .b(EX530), .O(N734) );
xor2 gate182( .a(N45), .b(N703), .O(N735) );
xor2 gate183( .a(N49), .b(N704), .O(N736) );
xor2 gate184( .a(N53), .b(N705), .O(N737) );
xor2 gate185( .a(N57), .b(N706), .O(N738) );
inv1 gate( .a(N61),.O(N61_NOT) );
inv1 gate( .a(N707),.O(N707_NOT));
and2 gate( .a(N61_NOT), .b(p213), .O(EX531) );
and2 gate( .a(N707_NOT), .b(EX531), .O(EX532) );
and2 gate( .a(N61), .b(p214), .O(EX533) );
and2 gate( .a(N707_NOT), .b(EX533), .O(EX534) );
and2 gate( .a(N61_NOT), .b(p215), .O(EX535) );
and2 gate( .a(N707), .b(EX535), .O(EX536) );
and2 gate( .a(N61), .b(p216), .O(EX537) );
and2 gate( .a(N707), .b(EX537), .O(EX538) );
or2  gate( .a(EX532), .b(EX534), .O(EX539) );
or2  gate( .a(EX536), .b(EX539), .O(EX540) );
or2  gate( .a(EX538), .b(EX540), .O(N739) );
inv1 gate( .a(N65),.O(N65_NOT) );
inv1 gate( .a(N708),.O(N708_NOT));
and2 gate( .a(N65_NOT), .b(p217), .O(EX541) );
and2 gate( .a(N708_NOT), .b(EX541), .O(EX542) );
and2 gate( .a(N65), .b(p218), .O(EX543) );
and2 gate( .a(N708_NOT), .b(EX543), .O(EX544) );
and2 gate( .a(N65_NOT), .b(p219), .O(EX545) );
and2 gate( .a(N708), .b(EX545), .O(EX546) );
and2 gate( .a(N65), .b(p220), .O(EX547) );
and2 gate( .a(N708), .b(EX547), .O(EX548) );
or2  gate( .a(EX542), .b(EX544), .O(EX549) );
or2  gate( .a(EX546), .b(EX549), .O(EX550) );
or2  gate( .a(EX548), .b(EX550), .O(N740) );
inv1 gate( .a(N69),.O(N69_NOT) );
inv1 gate( .a(N709),.O(N709_NOT));
and2 gate( .a(N69_NOT), .b(p221), .O(EX551) );
and2 gate( .a(N709_NOT), .b(EX551), .O(EX552) );
and2 gate( .a(N69), .b(p222), .O(EX553) );
and2 gate( .a(N709_NOT), .b(EX553), .O(EX554) );
and2 gate( .a(N69_NOT), .b(p223), .O(EX555) );
and2 gate( .a(N709), .b(EX555), .O(EX556) );
and2 gate( .a(N69), .b(p224), .O(EX557) );
and2 gate( .a(N709), .b(EX557), .O(EX558) );
or2  gate( .a(EX552), .b(EX554), .O(EX559) );
or2  gate( .a(EX556), .b(EX559), .O(EX560) );
or2  gate( .a(EX558), .b(EX560), .O(N741) );
xor2 gate189( .a(N73), .b(N710), .O(N742) );
inv1 gate( .a(N77),.O(N77_NOT) );
inv1 gate( .a(N711),.O(N711_NOT));
and2 gate( .a(N77_NOT), .b(p225), .O(EX561) );
and2 gate( .a(N711_NOT), .b(EX561), .O(EX562) );
and2 gate( .a(N77), .b(p226), .O(EX563) );
and2 gate( .a(N711_NOT), .b(EX563), .O(EX564) );
and2 gate( .a(N77_NOT), .b(p227), .O(EX565) );
and2 gate( .a(N711), .b(EX565), .O(EX566) );
and2 gate( .a(N77), .b(p228), .O(EX567) );
and2 gate( .a(N711), .b(EX567), .O(EX568) );
or2  gate( .a(EX562), .b(EX564), .O(EX569) );
or2  gate( .a(EX566), .b(EX569), .O(EX570) );
or2  gate( .a(EX568), .b(EX570), .O(N743) );
xor2 gate191( .a(N81), .b(N712), .O(N744) );
xor2 gate192( .a(N85), .b(N713), .O(N745) );
inv1 gate( .a(N89),.O(N89_NOT) );
inv1 gate( .a(N714),.O(N714_NOT));
and2 gate( .a(N89_NOT), .b(p229), .O(EX571) );
and2 gate( .a(N714_NOT), .b(EX571), .O(EX572) );
and2 gate( .a(N89), .b(p230), .O(EX573) );
and2 gate( .a(N714_NOT), .b(EX573), .O(EX574) );
and2 gate( .a(N89_NOT), .b(p231), .O(EX575) );
and2 gate( .a(N714), .b(EX575), .O(EX576) );
and2 gate( .a(N89), .b(p232), .O(EX577) );
and2 gate( .a(N714), .b(EX577), .O(EX578) );
or2  gate( .a(EX572), .b(EX574), .O(EX579) );
or2  gate( .a(EX576), .b(EX579), .O(EX580) );
or2  gate( .a(EX578), .b(EX580), .O(N746) );
inv1 gate( .a(N93),.O(N93_NOT) );
inv1 gate( .a(N715),.O(N715_NOT));
and2 gate( .a(N93_NOT), .b(p233), .O(EX581) );
and2 gate( .a(N715_NOT), .b(EX581), .O(EX582) );
and2 gate( .a(N93), .b(p234), .O(EX583) );
and2 gate( .a(N715_NOT), .b(EX583), .O(EX584) );
and2 gate( .a(N93_NOT), .b(p235), .O(EX585) );
and2 gate( .a(N715), .b(EX585), .O(EX586) );
and2 gate( .a(N93), .b(p236), .O(EX587) );
and2 gate( .a(N715), .b(EX587), .O(EX588) );
or2  gate( .a(EX582), .b(EX584), .O(EX589) );
or2  gate( .a(EX586), .b(EX589), .O(EX590) );
or2  gate( .a(EX588), .b(EX590), .O(N747) );
inv1 gate( .a(N97),.O(N97_NOT) );
inv1 gate( .a(N716),.O(N716_NOT));
and2 gate( .a(N97_NOT), .b(p237), .O(EX591) );
and2 gate( .a(N716_NOT), .b(EX591), .O(EX592) );
and2 gate( .a(N97), .b(p238), .O(EX593) );
and2 gate( .a(N716_NOT), .b(EX593), .O(EX594) );
and2 gate( .a(N97_NOT), .b(p239), .O(EX595) );
and2 gate( .a(N716), .b(EX595), .O(EX596) );
and2 gate( .a(N97), .b(p240), .O(EX597) );
and2 gate( .a(N716), .b(EX597), .O(EX598) );
or2  gate( .a(EX592), .b(EX594), .O(EX599) );
or2  gate( .a(EX596), .b(EX599), .O(EX600) );
or2  gate( .a(EX598), .b(EX600), .O(N748) );
xor2 gate196( .a(N101), .b(N717), .O(N749) );
xor2 gate197( .a(N105), .b(N718), .O(N750) );
inv1 gate( .a(N109),.O(N109_NOT) );
inv1 gate( .a(N719),.O(N719_NOT));
and2 gate( .a(N109_NOT), .b(p241), .O(EX601) );
and2 gate( .a(N719_NOT), .b(EX601), .O(EX602) );
and2 gate( .a(N109), .b(p242), .O(EX603) );
and2 gate( .a(N719_NOT), .b(EX603), .O(EX604) );
and2 gate( .a(N109_NOT), .b(p243), .O(EX605) );
and2 gate( .a(N719), .b(EX605), .O(EX606) );
and2 gate( .a(N109), .b(p244), .O(EX607) );
and2 gate( .a(N719), .b(EX607), .O(EX608) );
or2  gate( .a(EX602), .b(EX604), .O(EX609) );
or2  gate( .a(EX606), .b(EX609), .O(EX610) );
or2  gate( .a(EX608), .b(EX610), .O(N751) );
inv1 gate( .a(N113),.O(N113_NOT) );
inv1 gate( .a(N720),.O(N720_NOT));
and2 gate( .a(N113_NOT), .b(p245), .O(EX611) );
and2 gate( .a(N720_NOT), .b(EX611), .O(EX612) );
and2 gate( .a(N113), .b(p246), .O(EX613) );
and2 gate( .a(N720_NOT), .b(EX613), .O(EX614) );
and2 gate( .a(N113_NOT), .b(p247), .O(EX615) );
and2 gate( .a(N720), .b(EX615), .O(EX616) );
and2 gate( .a(N113), .b(p248), .O(EX617) );
and2 gate( .a(N720), .b(EX617), .O(EX618) );
or2  gate( .a(EX612), .b(EX614), .O(EX619) );
or2  gate( .a(EX616), .b(EX619), .O(EX620) );
or2  gate( .a(EX618), .b(EX620), .O(N752) );
inv1 gate( .a(N117),.O(N117_NOT) );
inv1 gate( .a(N721),.O(N721_NOT));
and2 gate( .a(N117_NOT), .b(p249), .O(EX621) );
and2 gate( .a(N721_NOT), .b(EX621), .O(EX622) );
and2 gate( .a(N117), .b(p250), .O(EX623) );
and2 gate( .a(N721_NOT), .b(EX623), .O(EX624) );
and2 gate( .a(N117_NOT), .b(p251), .O(EX625) );
and2 gate( .a(N721), .b(EX625), .O(EX626) );
and2 gate( .a(N117), .b(p252), .O(EX627) );
and2 gate( .a(N721), .b(EX627), .O(EX628) );
or2  gate( .a(EX622), .b(EX624), .O(EX629) );
or2  gate( .a(EX626), .b(EX629), .O(EX630) );
or2  gate( .a(EX628), .b(EX630), .O(N753) );
inv1 gate( .a(N121),.O(N121_NOT) );
inv1 gate( .a(N722),.O(N722_NOT));
and2 gate( .a(N121_NOT), .b(p253), .O(EX631) );
and2 gate( .a(N722_NOT), .b(EX631), .O(EX632) );
and2 gate( .a(N121), .b(p254), .O(EX633) );
and2 gate( .a(N722_NOT), .b(EX633), .O(EX634) );
and2 gate( .a(N121_NOT), .b(p255), .O(EX635) );
and2 gate( .a(N722), .b(EX635), .O(EX636) );
and2 gate( .a(N121), .b(p256), .O(EX637) );
and2 gate( .a(N722), .b(EX637), .O(EX638) );
or2  gate( .a(EX632), .b(EX634), .O(EX639) );
or2  gate( .a(EX636), .b(EX639), .O(EX640) );
or2  gate( .a(EX638), .b(EX640), .O(N754) );
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule
