
module c3540 (N1,N13,N20,N33,N41,N45,N50,N58,N68,N77,
              N87,N97,N107,N116,N124,N125,N128,N132,N137,N143,
              N150,N159,N169,N179,N190,N200,N213,N222,N223,N226,
              N232,N238,N244,N250,N257,N264,N270,N274,N283,N294,
              N303,N311,N317,N322,N326,N329,N330,N343,N349,N350,
              N1713,N1947,N3195,N3833,N3987,N4028,N4145,N4589,N4667,N4815,
              N4944,N5002,N5045,N5047,N5078,N5102,N5120,N5121,N5192,N5231,
              N5360,N5361);

input N1_new,N13_new,N20_new,N33_new,N41_new,N45_new,N50_new,N58_new,N68_new,N77_new,
      N87_new,N97_new,N107_new,N116_new,N124_new,N125_new,N128_new,N132_new,N137_new,N143_new,
      N150_new,N159_new,N169_new,N179_new,N190_new,N200_new,N213_new,N222_new,N223_new,N226_new,
      N232_new,N238_new,N244_new,N250_new,N257_new,N264_new,N270_new,N274_new,N283_new,N294_new,
      N303_new,N311_new,N317_new,N322_new,N326_new,N329_new,N330_new,N343_new,N349_new,N350_new;

input p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,
        p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,
        p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,
        p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,
        p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,
        p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,
        p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,
        p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,
        p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,
        p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,
        p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,
        p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,
        p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,
        p131,p132,p133,p134,p135,p136,p137,p138,p139,p140,
        p141,p142,p143,p144,p145,p146,p147,p148,p149,p150,
        p151,p152,p153,p154,p155,p156,p157,p158,p159,p160,
        p161,p162,p163,p164,p165,p166,p167,p168,p169,p170,
        p171,p172,p173,p174,p175,p176,p177,p178,p179,p180,
        p181,p182,p183,p184,p185,p186,p187,p188,p189,p190,
        p191,p192,p193,p194,p195,p196,p197,p198,p199,p200,
        p201,p202,p203,p204,p205,p206,p207,p208,p209,p210,
        p211,p212,p213,p214,p215,p216,p217,p218,p219,p220,
        p221,p222,p223,p224,p225,p226,p227,p228,p229,p230,
        p231,p232,p233,p234,p235,p236,p237,p238,p239,p240,
        p241,p242,p243,p244,p245,p246,p247,p248,p249,p250,
        p251,p252,p253,p254,p255,p256,p257,p258,p259,p260,
        p261,p262,p263,p264,p265,p266,p267,p268,p269,p270,
        p271,p272,p273,p274,p275,p276,p277,p278,p279,p280,
        p281,p282,p283,p284,p285,p286,p287,p288,p289,p290,
        p291,p292,p293,p294,p295,p296,p297,p298,p299,p300,
        p301,p302,p303,p304,p305,p306,p307,p308,p309,p310,
        p311,p312,p313,p314,p315,p316,p317,p318,p319,p320,
        p321,p322,p323,p324,p325,p326,p327,p328,p329,p330,
        p331,p332,p333,p334,p335,p336,p337,p338,p339,p340,
        p341,p342,p343,p344,p345,p346,p347,p348,p349,p350,
        p351,p352,p353,p354,p355,p356,p357,p358,p359,p360,
        p361,p362,p363,p364,p365,p366,p367,p368,p369,p370,
        p371,p372,p373,p374,p375,p376,p377,p378,p379,p380,
        p381,p382,p383,p384,p385,p386,p387,p388,p389,p390,
        p391,p392,p393,p394,p395,p396,p397,p398,p399,p400,
        p401,p402,p403,p404,p405,p406,p407,p408,p409,p410,
        p411,p412,p413,p414,p415,p416,p417,p418,p419,p420,
        p421,p422,p423,p424,p425,p426,p427,p428,p429,p430,
        p431,p432,p433,p434,p435,p436,p437,p438,p439,p440,
        p441,p442,p443,p444,p445,p446,p447,p448,p449,p450,
        p451,p452,p453,p454,p455,p456,p457,p458,p459,p460,
        p461,p462,p463,p464,p465,p466,p467,p468,p469,p470,
        p471,p472,p473,p474,p475,p476,p477,p478,p479,p480,
        p481,p482,p483,p484,p485,p486,p487,p488,p489,p490,
        p491,p492,p493,p494,p495,p496,p497,p498,p499,p500,
        p501,p502,p503,p504,p505,p506,p507,p508,p509,p510,
        p511,p512,p513,p514,p515,p516,p517,p518,p519,p520,
        p521,p522,p523,p524,p525,p526,p527,p528,p529,p530,
        p531,p532,p533,p534,p535,p536,p537,p538,p539,p540,
        p541,p542,p543,p544,p545,p546,p547,p548,p549,p550,
        p551,p552,p553,p554,p555,p556,p557,p558,p559,p560,
        p561,p562,p563,p564,p565,p566,p567,p568,p569,p570,
        p571,p572,p573,p574,p575,p576,p577,p578,p579,p580,
        p581,p582,p583,p584,p585,p586,p587,p588,p589,p590,
        p591,p592,p593,p594,p595,p596,p597,p598,p599,p600,
        p601,p602,p603,p604,p605,p606,p607,p608,p609,p610,
        p611,p612,p613,p614,p615,p616,p617,p618,p619,p620,
        p621,p622,p623,p624,p625,p626,p627,p628,p629,p630,
        p631,p632,p633,p634,p635,p636,p637,p638,p639,p640,
        p641,p642,p643,p644,p645,p646,p647,p648,p649,p650,
        p651,p652,p653,p654,p655,p656,X_1,X_2,X_3,X_4,X_5,X_6,X_7,X_8,X_9,X_10,X_11,X_12,X_13,X_14,X_15,X_16,X_17,X_18,X_19,X_20,X_21,X_22,X_23,X_24,X_25,X_26,X_27,X_28,X_29,X_30,X_31,X_32,X_33,X_34,X_35,X_36,X_37,X_38,X_39,X_40,X_41,X_42,X_43,X_44,X_45,X_46,X_47,X_48,X_49,X_50,X_51,X_52,X_53,X_54,X_55,X_56,X_57,X_58,X_59,X_60,X_61,X_62,X_63,X_64,X_65,X_66,X_67,X_68,X_69,X_70,X_71,X_72;

output N1713_new,N1947_new,N3195_new,N3833_new,N3987_new,N4028_new,N4145_new,N4589_new,N4667_new,N4815_new,
       N4944_new,N5002_new,N5045_new,N5047_new,N5078_new,N5102_new,N5120_new,N5121_new,N5192_new,N5231_new,
       N5360_new,N5361_new;

wire N655,N665,N670,N679,N683,N686,N690,N699,N702,N706,
     N715,N724,N727,N736,N740,N749,N753,N763,N768,N769,
     N772,N779,N782,N786,N793,N794,N798,N803,N820,N821,
     N825,N829,N832,N835,N836,N839,N842,N845,N848,N851,
     N854,N858,N861,N864,N867,N870,N874,N877,N880,N883,
     N886,N889,N890,N891,N892,N895,N896,N913,N914,N915,
     N916,N917,N920,N923,N926,N929,N932,N935,N938,N941,
     N944,N947,N950,N953,N956,N959,N962,N965,N1067,N1117,
     N1179,N1196,N1197,N1202,N1219,N1250,N1251,N1252,N1253,N1254,
     N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,
     N1267,N1268,N1271,N1272,N1273,N1276,N1279,N1298,N1302,N1306,
     N1315,N1322,N1325,N1328,N1331,N1334,N1337,N1338,N1339,N1340,
     N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,
     N1353,N1358,N1363,N1366,N1369,N1384,N1401,N1402,N1403,N1404,
     N1405,N1406,N1407,N1408,N1409,N1426,N1427,N1452,N1459,N1460,
     N1461,N1464,N1467,N1468,N1469,N1470,N1471,N1474,N1475,N1478,
     N1481,N1484,N1487,N1490,N1493,N1496,N1499,N1502,N1505,N1507,
     N1508,N1509,N1510,N1511,N1512,N1520,N1562,N1579,N1580,N1581,
     N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,
     N1592,N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1643,
     N1644,N1645,N1646,N1647,N1648,N1649,N1650,N1667,N1670,N1673,
     N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1691,N1692,N1693,
     N1694,N1714,N1715,N1718,N1721,N1722,N1725,N1726,N1727,N1728,
     N1729,N1730,N1731,N1735,N1736,N1737,N1738,N1747,N1756,N1761,
     N1764,N1765,N1766,N1767,N1768,N1769,N1770,N1787,N1788,N1789,
     N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,N1798,N1799,
     N1800,N1801,N1802,N1803,N1806,N1809,N1812,N1815,N1818,N1821,
     N1824,N1833,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,
     N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,
     N1860,N1861,N1862,N1863,N1864,N1869,N1870,N1873,N1874,N1875,
     N1878,N1879,N1880,N1883,N1884,N1885,N1888,N1889,N1890,N1893,
     N1894,N1895,N1898,N1899,N1900,N1903,N1904,N1905,N1908,N1909,
     N1912,N1913,N1917,N1922,N1926,N1930,N1933,N1936,N1939,N1940,
     N1941,N1942,N1943,N1944,N1945,N1946,N1960,N1961,N1966,N1981,
     N1982,N1983,N1986,N1987,N1988,N1989,N1990,N1991,N2022,N2023,
     N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,
     N2034,N2035,N2036,N2037,N2038,N2043,N2052,N2057,N2068,N2073,
     N2078,N2083,N2088,N2093,N2098,N2103,N2121,N2122,N2123,N2124,
     N2125,N2126,N2127,N2128,N2133,N2134,N2135,N2136,N2137,N2138,
     N2139,N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,N2149,
     N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,N2158,N2175,
     N2178,N2179,N2180,N2181,N2183,N2184,N2185,N2188,N2191,N2194,
     N2197,N2200,N2203,N2206,N2209,N2210,N2211,N2212,N2221,N2230,
     N2231,N2232,N2233,N2234,N2235,N2236,N2237,N2238,N2239,N2240,
     N2241,N2242,N2243,N2244,N2245,N2270,N2277,N2282,N2287,N2294,
     N2299,N2304,N2307,N2310,N2313,N2316,N2319,N2322,N2325,N2328,
     N2331,N2334,N2341,N2342,N2347,N2348,N2349,N2350,N2351,N2352,
     N2353,N2354,N2355,N2374,N2375,N2376,N2379,N2398,N2417,N2418,
     N2419,N2420,N2421,N2422,N2425,N2426,N2427,N2430,N2431,N2432,
     N2435,N2436,N2437,N2438,N2439,N2440,N2443,N2444,N2445,N2448,
     N2449,N2450,N2467,N2468,N2469,N2470,N2471,N2474,N2475,N2476,
     N2477,N2478,N2481,N2482,N2483,N2486,N2487,N2488,N2497,N2506,
     N2515,N2524,N2533,N2542,N2551,N2560,N2569,N2578,N2587,N2596,
     N2605,N2614,N2623,N2632,N2633,N2634,N2635,N2636,N2637,N2638,
     N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,N2647,N2648,
     N2652,N2656,N2659,N2662,N2666,N2670,N2673,N2677,N2681,N2684,
     N2688,N2692,N2697,N2702,N2706,N2710,N2715,N2719,N2723,N2728,
     N2729,N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,
     N2739,N2740,N2741,N2742,N2743,N2744,N2745,N2746,N2748,N2749,
     N2750,N2751,N2754,N2755,N2756,N2757,N2758,N2761,N2764,N2768,
     N2769,N2898,N2899,N2900,N2901,N2962,N2966,N2967,N2970,N2973,
     N2977,N2980,N2984,N2985,N2986,N2987,N2988,N2989,N2990,N2991,
     N2992,N2993,N2994,N2995,N2996,N2997,N2998,N2999,N3000,N3001,
     N3002,N3003,N3004,N3005,N3006,N3007,N3008,N3009,N3010,N3011,
     N3012,N3013,N3014,N3015,N3016,N3017,N3018,N3019,N3020,N3021,
     N3022,N3023,N3024,N3025,N3026,N3027,N3028,N3029,N3030,N3031,
     N3032,N3033,N3034,N3035,N3036,N3037,N3038,N3039,N3040,N3041,
     N3042,N3043,N3044,N3045,N3046,N3047,N3048,N3049,N3050,N3051,
     N3052,N3053,N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061,
     N3062,N3063,N3064,N3065,N3066,N3067,N3068,N3069,N3070,N3071,
     N3072,N3073,N3074,N3075,N3076,N3077,N3078,N3079,N3080,N3081,
     N3082,N3083,N3084,N3085,N3086,N3087,N3088,N3089,N3090,N3091,
     N3092,N3093,N3094,N3095,N3096,N3097,N3098,N3099,N3100,N3101,
     N3102,N3103,N3104,N3105,N3106,N3107,N3108,N3109,N3110,N3111,
     N3112,N3115,N3118,N3119,N3122,N3125,N3128,N3131,N3134,N3135,
     N3138,N3141,N3142,N3145,N3148,N3149,N3152,N3155,N3158,N3161,
     N3164,N3165,N3168,N3171,N3172,N3175,N3178,N3181,N3184,N3187,
     N3190,N3191,N3192,N3193,N3194,N3196,N3206,N3207,N3208,N3209,
     N3210,N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,N3219,
     N3220,N3221,N3222,N3223,N3224,N3225,N3226,N3227,N3228,N3229,
     N3230,N3231,N3232,N3233,N3234,N3235,N3236,N3237,N3238,N3239,
     N3240,N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3248,N3249,
     N3250,N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,N3259,
     N3260,N3261,N3262,N3263,N3264,N3265,N3266,N3267,N3268,N3269,
     N3270,N3271,N3272,N3273,N3274,N3275,N3276,N3277,N3278,N3279,
     N3280,N3281,N3282,N3283,N3284,N3285,N3286,N3287,N3288,N3289,
     N3290,N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,N3299,
     N3300,N3301,N3302,N3303,N3304,N3305,N3306,N3307,N3308,N3309,
     N3310,N3311,N3312,N3313,N3314,N3315,N3316,N3317,N3318,N3319,
     N3320,N3321,N3322,N3323,N3324,N3325,N3326,N3327,N3328,N3329,
     N3330,N3331,N3332,N3333,N3334,N3383,N3384,N3387,N3388,N3389,
     N3390,N3391,N3392,N3393,N3394,N3395,N3396,N3397,N3398,N3399,
     N3400,N3401,N3402,N3403,N3404,N3405,N3406,N3407,N3410,N3413,
     N3414,N3415,N3419,N3423,N3426,N3429,N3430,N3431,N3434,N3437,
     N3438,N3439,N3442,N3445,N3446,N3447,N3451,N3455,N3458,N3461,
     N3462,N3463,N3466,N3469,N3470,N3471,N3472,N3475,N3478,N3481,
     N3484,N3487,N3490,N3493,N3496,N3499,N3502,N3505,N3508,N3511,
     N3514,N3517,N3520,N3523,N3534,N3535,N3536,N3537,N3538,N3539,
     N3540,N3541,N3542,N3543,N3544,N3545,N3546,N3547,N3548,N3549,
     N3550,N3551,N3552,N3557,N3568,N3573,N3578,N3589,N3594,N3605,
     N3626,N3627,N3628,N3629,N3630,N3631,N3632,N3633,N3634,N3635,
     N3636,N3637,N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,
     N3648,N3651,N3652,N3653,N3654,N3657,N3658,N3661,N3662,N3663,
     N3664,N3667,N3670,N3671,N3672,N3673,N3676,N3677,N3680,N3681,
     N3682,N3685,N3686,N3687,N3688,N3689,N3690,N3693,N3694,N3695,
     N3696,N3697,N3700,N3703,N3704,N3705,N3706,N3707,N3708,N3711,
     N3712,N3713,N3714,N3715,N3716,N3717,N3718,N3719,N3720,N3721,
     N3731,N3734,N3740,N3743,N3753,N3756,N3762,N3765,N3766,N3773,
     N3774,N3775,N3776,N3777,N3778,N3779,N3780,N3786,N3789,N3800,
     N3803,N3809,N3812,N3815,N3818,N3821,N3824,N3827,N3830,N3834,
     N3835,N3838,N3845,N3850,N3855,N3858,N3861,N3865,N3868,N3884,
     N3885,N3894,N3895,N3898,N3899,N3906,N3911,N3912,N3913,N3916,
     N3917,N3920,N3921,N3924,N3925,N3926,N3930,N3931,N3932,N3935,
     N3936,N3937,N3940,N3947,N3948,N3950,N3953,N3956,N3959,N3962,
     N3965,N3968,N3971,N3974,N3977,N3980,N3983,N3992,N3996,N4013,
     N4029,N4030,N4031,N4032,N4033,N4034,N4035,N4042,N4043,N4044,
     N4045,N4046,N4047,N4048,N4049,N4050,N4051,N4052,N4053,N4054,
     N4055,N4056,N4057,N4058,N4059,N4062,N4065,N4066,N4067,N4070,
     N4073,N4074,N4075,N4076,N4077,N4078,N4079,N4080,N4085,N4086,
     N4088,N4090,N4091,N4094,N4098,N4101,N4104,N4105,N4106,N4107,
     N4108,N4109,N4110,N4111,N4112,N4113,N4114,N4115,N4116,N4119,
     N4122,N4123,N4126,N4127,N4128,N4139,N4142,N4146,N4147,N4148,
     N4149,N4150,N4151,N4152,N4153,N4154,N4161,N4167,N4174,N4182,
     N4186,N4189,N4190,N4191,N4192,N4193,N4194,N4195,N4196,N4197,
     N4200,N4203,N4209,N4213,N4218,N4223,N4238,N4239,N4241,N4242,
     N4247,N4251,N4252,N4253,N4254,N4255,N4256,N4257,N4258,N4283,
     N4284,N4287,N4291,N4295,N4296,N4299,N4303,N4304,N4305,N4310,
     N4316,N4317,N4318,N4319,N4322,N4325,N4326,N4327,N4328,N4329,
     N4330,N4331,N4335,N4338,N4341,N4344,N4347,N4350,N4353,N4356,
     N4359,N4362,N4365,N4368,N4371,N4376,N4377,N4387,N4390,N4393,
     N4398,N4413,N4416,N4421,N4427,N4430,N4435,N4442,N4443,N4446,
     N4447,N4448,N4452,N4458,N4461,N4462,N4463,N4464,N4465,N4468,
     N4472,N4475,N4479,N4484,N4486,N4487,N4491,N4493,N4496,N4497,
     N4498,N4503,N4506,N4507,N4508,N4509,N4510,N4511,N4515,N4526,
     N4527,N4528,N4529,N4530,N4531,N4534,N4537,N4540,N4545,N4549,
     N4552,N4555,N4558,N4559,N4562,N4563,N4564,N4568,N4569,N4572,
     N4573,N4576,N4581,N4584,N4587,N4588,N4593,N4596,N4597,N4599,
     N4602,N4603,N4608,N4613,N4616,N4619,N4623,N4628,N4629,N4630,
     N4635,N4636,N4640,N4641,N4642,N4643,N4644,N4647,N4650,N4656,
     N4659,N4664,N4668,N4669,N4670,N4673,N4674,N4675,N4676,N4677,
     N4678,N4679,N4687,N4688,N4691,N4694,N4697,N4700,N4704,N4705,
     N4706,N4707,N4708,N4711,N4716,N4717,N4721,N4722,N4726,N4727,
     N4730,N4733,N4740,N4743,N4747,N4748,N4749,N4750,N4753,N4754,
     N4755,N4756,N4757,N4769,N4772,N4775,N4778,N4786,N4787,N4788,
     N4789,N4794,N4797,N4800,N4805,N4808,N4812,N4816,N4817,N4818,
     N4822,N4823,N4826,N4829,N4830,N4831,N4838,N4844,N4847,N4850,
     N4854,N4859,N4860,N4868,N4870,N4872,N4873,N4876,N4880,N4885,
     N4889,N4895,N4896,N4897,N4898,N4899,N4900,N4901,N4902,N4904,
     N4905,N4906,N4907,N4913,N4916,N4920,N4921,N4924,N4925,N4926,
     N4928,N4929,N4930,N4931,N4937,N4940,N4946,N4949,N4950,N4951,
     N4952,N4953,N4954,N4957,N4964,N4965,N4968,N4969,N4970,N4973,
     N4978,N4979,N4980,N4981,N4982,N4983,N4984,N4985,N4988,N4991,
     N4996,N4999,N5007,N5010,N5013,N5018,N5021,N5026,N5029,N5030,
     N5039,N5042,N5046,N5050,N5055,N5058,N5061,N5066,N5070,N5080,
     N5085,N5094,N5095,N5097,N5103,N5108,N5109,N5110,N5111,N5114,
     N5117,N5122,N5125,N5128,N5133,N5136,N5139,N5145,N5151,N5154,
     N5159,N5160,N5163,N5166,N5173,N5174,N5177,N5182,N5183,N5184,
     N5188,N5193,N5196,N5197,N5198,N5199,N5201,N5203,N5205,N5209,
     N5212,N5215,N5217,N5219,N5220,N5221,N5222,N5223,N5224,N5225,
     N5228,N5232,N5233,N5234,N5235,N5236,N5240,N5242,N5243,N5245,
     N5246,N5250,N5253,N5254,N5257,N5258,N5261,N5266,N5269,N5277,
     N5278,N5279,N5283,N5284,N5285,N5286,N5289,N5292,N5295,N5298,
     N5303,N5306,N5309,N5312,N5313,N5322,N5323,N5324,N5327,N5332,
     N5335,N5340,N5341,N5344,N5345,N5348,N5349,N5350,N5351,N5352,
     N5353,N5354,N5355,N5356,N5357,N5358,N5359,
     N257_NOT,N264_NOT,N13_NOT,N20_NOT,N33_NOT,N41_NOT,N41_NOT,N45_NOT,N20_NOT,N200_NOT,
     N20_NOT,N200_NOT,N349_NOT,N33_NOT,N895_NOT,N169_NOT,N915_NOT,N1_NOT,N916_NOT,N1_NOT,
     N226_NOT,N655_NOT,N232_NOT,N670_NOT,N250_NOT,N715_NOT,N257_NOT,N727_NOT,N264_NOT,N740_NOT,
     N920_NOT,N923_NOT,N920_NOT,N923_NOT,N702_NOT,N1250_NOT,N77_NOT,N1348_NOT,N803_NOT,N1117_NOT,
     N238_NOT,N1405_NOT,N244_NOT,N1406_NOT,N257_NOT,N1408_NOT,N1502_NOT,N1344_NOT,N150_NOT,N1580_NOT,
     N851_NOT,N1582_NOT,N858_NOT,N1587_NOT,N891_NOT,N1366_NOT,N786_NOT,N1298_NOT,N68_NOT,N1409_NOT,
     N1202_NOT,N1409_NOT,N1202_NOT,N1409_NOT,N1693_NOT,N1694_NOT,N223_NOT,N1850_NOT,N107_NOT,N1855_NOT,
     N303_NOT,N1863_NOT,N950_NOT,N1939_NOT,N1481_NOT,N1944_NOT,N1487_NOT,N1946_NOT,N1353_NOT,N1812_NOT,
     N1930_NOT,N350_NOT,N1930_NOT,N350_NOT,N1933_NOT,N2142_NOT,N763_NOT,N2154_NOT,N1725_NOT,N2156_NOT,
     N1520_NOT,N2180_NOT,N1721_NOT,N2181_NOT,N2052_NOT,N2238_NOT,N2052_NOT,N2239_NOT,N2038_NOT,N2242_NOT,
     N2348_NOT,N1729_NOT,N2175_NOT,N1334_NOT,N2349_NOT,N2183_NOT,N2212_NOT,N1833_NOT,N1562_NOT,N2158_NOT,
     N1562_NOT,N2158_NOT,N2316_NOT,N2467_NOT,N2325_NOT,N2475_NOT,N1520_NOT,N2481_NOT,N1722_NOT,N2482_NOT,
     N665_NOT,N2633_NOT,N2768_NOT,N1674_NOT,N1913_NOT,N2673_NOT,N1922_NOT,N2715_NOT,N159_NOT,N2985_NOT,
     N150_NOT,N2986_NOT,N143_NOT,N2987_NOT,N132_NOT,N2989_NOT,N159_NOT,N2994_NOT,N655_NOT,N3020_NOT,
     N715_NOT,N3025_NOT,N670_NOT,N3028_NOT,N150_NOT,N3032_NOT,N690_NOT,N3036_NOT,N283_NOT,N3048_NOT,
     N727_NOT,N3053_NOT,N753_NOT,N3062_NOT,N283_NOT,N3063_NOT,N715_NOT,N3066_NOT,N740_NOT,N3068_NOT,
     N311_NOT,N3072_NOT,N715_NOT,N3073_NOT,N727_NOT,N3074_NOT,N740_NOT,N3075_NOT,N317_NOT,N3080_NOT,
     N283_NOT,N3084_NOT,N294_NOT,N3085_NOT,N753_NOT,N3090_NOT,N283_NOT,N3091_NOT,N303_NOT,N3093_NOT,
     N317_NOT,N3095_NOT,N283_NOT,N3098_NOT,N329_NOT,N3104_NOT,N3196_NOT,N1736_NOT,N3387_NOT,N2350_NOT,
     N3392_NOT,N1843_NOT,N3396_NOT,N1847_NOT,N3407_NOT,N3410_NOT,N3439_NOT,N3442_NOT,N3475_NOT,N3630_NOT,
     N3481_NOT,N3626_NOT,N3478_NOT,N3627_NOT,N3636_NOT,N2636_NOT,N3637_NOT,N2638_NOT,N3641_NOT,N2646_NOT,
     N3705_NOT,N3706_NOT,N3707_NOT,N3708_NOT,N3700_NOT,N3628_NOT,N3677_NOT,N1926_NOT,N3487_NOT,N3776_NOT,
     N3956_NOT,N3685_NOT,N3980_NOT,N3694_NOT,N3508_NOT,N4065_NOT,N4073_NOT,N4074_NOT,N4075_NOT,N4029_NOT,
     N4079_NOT,N4033_NOT,N4090_NOT,N4055_NOT,N3824_NOT,N4115_NOT,N4148_NOT,N2232_NOT,N4161_NOT,N4127_NOT,
     N4174_NOT,N4035_NOT,N3992_NOT,N4283_NOT,N4251_NOT,N2730_NOT,N4253_NOT,N2734_NOT,N4254_NOT,N2736_NOT,
     N4255_NOT,N2738_NOT,N4258_NOT,N2744_NOT,N330_NOT,N4316_NOT,N4377_NOT,N2740_NOT,N4427_NOT,N4241_NOT,
     N965_NOT,N4464_NOT,N330_NOT,N4443_NOT,N4310_NOT,N4465_NOT,N4362_NOT,N4529_NOT,N4559_NOT,N2128_NOT,
     N4616_NOT,N4239_NOT,N4186_NOT,N4635_NOT,N4365_NOT,N4640_NOT,N4629_NOT,N4668_NOT,N4435_NOT,N4673_NOT,
     N4493_NOT,N4676_NOT,N4531_NOT,N4747_NOT,N4711_NOT,N2735_NOT,N4717_NOT,N4468_NOT,N4786_NOT,N4748_NOT,
     N4854_NOT,N4872_NOT,N4895_NOT,N2184_NOT,N4930_NOT,N4905_NOT,N4953_NOT,N2739_NOT,N4950_NOT,N4969_NOT,
     N4981_NOT,N4982_NOT,N5007_NOT,N2729_NOT,N5050_NOT,N5050_NOT,N1461_NOT,N5080_NOT,N213_NOT,N5193_NOT,
     N4937_NOT,N5197_NOT,N5205_NOT,N5217_NOT,N5198_NOT,N5221_NOT,N5232_NOT,N5245_NOT,N5295_NOT,N5284_NOT,
     N5324_NOT,N5323_NOT,N5327_NOT,N5322_NOT,N5306_NOT,N5344_NOT,N5349_NOT,N5355_NOT,EX1,EX2,EX3,EX4,EX5,EX6,EX7,EX8,EX9,EX10,
     EX11,EX12,EX13,EX14,EX15,EX16,EX17,EX18,EX19,EX20,
     EX21,EX22,EX23,EX24,EX25,EX26,EX27,EX28,EX29,EX30,
     EX31,EX32,EX33,EX34,EX35,EX36,EX37,EX38,EX39,EX40,
     EX41,EX42,EX43,EX44,EX45,EX46,EX47,EX48,EX49,EX50,
     EX51,EX52,EX53,EX54,EX55,EX56,EX57,EX58,EX59,EX60,
     EX61,EX62,EX63,EX64,EX65,EX66,EX67,EX68,EX69,EX70,
     EX71,EX72,EX73,EX74,EX75,EX76,EX77,EX78,EX79,EX80,
     EX81,EX82,EX83,EX84,EX85,EX86,EX87,EX88,EX89,EX90,
     EX91,EX92,EX93,EX94,EX95,EX96,EX97,EX98,EX99,EX100,
     EX101,EX102,EX103,EX104,EX105,EX106,EX107,EX108,EX109,EX110,
     EX111,EX112,EX113,EX114,EX115,EX116,EX117,EX118,EX119,EX120,
     EX121,EX122,EX123,EX124,EX125,EX126,EX127,EX128,EX129,EX130,
     EX131,EX132,EX133,EX134,EX135,EX136,EX137,EX138,EX139,EX140,
     EX141,EX142,EX143,EX144,EX145,EX146,EX147,EX148,EX149,EX150,
     EX151,EX152,EX153,EX154,EX155,EX156,EX157,EX158,EX159,EX160,
     EX161,EX162,EX163,EX164,EX165,EX166,EX167,EX168,EX169,EX170,
     EX171,EX172,EX173,EX174,EX175,EX176,EX177,EX178,EX179,EX180,
     EX181,EX182,EX183,EX184,EX185,EX186,EX187,EX188,EX189,EX190,
     EX191,EX192,EX193,EX194,EX195,EX196,EX197,EX198,EX199,EX200,
     EX201,EX202,EX203,EX204,EX205,EX206,EX207,EX208,EX209,EX210,
     EX211,EX212,EX213,EX214,EX215,EX216,EX217,EX218,EX219,EX220,
     EX221,EX222,EX223,EX224,EX225,EX226,EX227,EX228,EX229,EX230,
     EX231,EX232,EX233,EX234,EX235,EX236,EX237,EX238,EX239,EX240,
     EX241,EX242,EX243,EX244,EX245,EX246,EX247,EX248,EX249,EX250,
     EX251,EX252,EX253,EX254,EX255,EX256,EX257,EX258,EX259,EX260,
     EX261,EX262,EX263,EX264,EX265,EX266,EX267,EX268,EX269,EX270,
     EX271,EX272,EX273,EX274,EX275,EX276,EX277,EX278,EX279,EX280,
     EX281,EX282,EX283,EX284,EX285,EX286,EX287,EX288,EX289,EX290,
     EX291,EX292,EX293,EX294,EX295,EX296,EX297,EX298,EX299,EX300,
     EX301,EX302,EX303,EX304,EX305,EX306,EX307,EX308,EX309,EX310,
     EX311,EX312,EX313,EX314,EX315,EX316,EX317,EX318,EX319,EX320,
     EX321,EX322,EX323,EX324,EX325,EX326,EX327,EX328,EX329,EX330,
     EX331,EX332,EX333,EX334,EX335,EX336,EX337,EX338,EX339,EX340,
     EX341,EX342,EX343,EX344,EX345,EX346,EX347,EX348,EX349,EX350,
     EX351,EX352,EX353,EX354,EX355,EX356,EX357,EX358,EX359,EX360,
     EX361,EX362,EX363,EX364,EX365,EX366,EX367,EX368,EX369,EX370,
     EX371,EX372,EX373,EX374,EX375,EX376,EX377,EX378,EX379,EX380,
     EX381,EX382,EX383,EX384,EX385,EX386,EX387,EX388,EX389,EX390,
     EX391,EX392,EX393,EX394,EX395,EX396,EX397,EX398,EX399,EX400,
     EX401,EX402,EX403,EX404,EX405,EX406,EX407,EX408,EX409,EX410,
     EX411,EX412,EX413,EX414,EX415,EX416,EX417,EX418,EX419,EX420,
     EX421,EX422,EX423,EX424,EX425,EX426,EX427,EX428,EX429,EX430,
     EX431,EX432,EX433,EX434,EX435,EX436,EX437,EX438,EX439,EX440,
     EX441,EX442,EX443,EX444,EX445,EX446,EX447,EX448,EX449,EX450,
     EX451,EX452,EX453,EX454,EX455,EX456,EX457,EX458,EX459,EX460,
     EX461,EX462,EX463,EX464,EX465,EX466,EX467,EX468,EX469,EX470,
     EX471,EX472,EX473,EX474,EX475,EX476,EX477,EX478,EX479,EX480,
     EX481,EX482,EX483,EX484,EX485,EX486,EX487,EX488,EX489,EX490,
     EX491,EX492,EX493,EX494,EX495,EX496,EX497,EX498,EX499,EX500,
     EX501,EX502,EX503,EX504,EX505,EX506,EX507,EX508,EX509,EX510,
     EX511,EX512,EX513,EX514,EX515,EX516,EX517,EX518,EX519,EX520,
     EX521,EX522,EX523,EX524,EX525,EX526,EX527,EX528,EX529,EX530,
     EX531,EX532,EX533,EX534,EX535,EX536,EX537,EX538,EX539,EX540,
     EX541,EX542,EX543,EX544,EX545,EX546,EX547,EX548,EX549,EX550,
     EX551,EX552,EX553,EX554,EX555,EX556,EX557,EX558,EX559,EX560,
     EX561,EX562,EX563,EX564,EX565,EX566,EX567,EX568,EX569,EX570,
     EX571,EX572,EX573,EX574,EX575,EX576,EX577,EX578,EX579,EX580,
     EX581,EX582,EX583,EX584,EX585,EX586,EX587,EX588,EX589,EX590,
     EX591,EX592,EX593,EX594,EX595,EX596,EX597,EX598,EX599,EX600,
     EX601,EX602,EX603,EX604,EX605,EX606,EX607,EX608,EX609,EX610,
     EX611,EX612,EX613,EX614,EX615,EX616,EX617,EX618,EX619,EX620,
     EX621,EX622,EX623,EX624,EX625,EX626,EX627,EX628,EX629,EX630,
     EX631,EX632,EX633,EX634,EX635,EX636,EX637,EX638,EX639,EX640,
     EX641,EX642,EX643,EX644,EX645,EX646,EX647,EX648,EX649,EX650,
     EX651,EX652,EX653,EX654,EX655,EX656,EX657,EX658,EX659,EX660,
     EX661,EX662,EX663,EX664,EX665,EX666,EX667,EX668,EX669,EX670,
     EX671,EX672,EX673,EX674,EX675,EX676,EX677,EX678,EX679,EX680,
     EX681,EX682,EX683,EX684,EX685,EX686,EX687,EX688,EX689,EX690,
     EX691,EX692,EX693,EX694,EX695,EX696,EX697,EX698,EX699,EX700,
     EX701,EX702,EX703,EX704,EX705,EX706,EX707,EX708,EX709,EX710,
     EX711,EX712,EX713,EX714,EX715,EX716,EX717,EX718,EX719,EX720,
     EX721,EX722,EX723,EX724,EX725,EX726,EX727,EX728,EX729,EX730,
     EX731,EX732,EX733,EX734,EX735,EX736,EX737,EX738,EX739,EX740,
     EX741,EX742,EX743,EX744,EX745,EX746,EX747,EX748,EX749,EX750,
     EX751,EX752,EX753,EX754,EX755,EX756,EX757,EX758,EX759,EX760,
     EX761,EX762,EX763,EX764,EX765,EX766,EX767,EX768,EX769,EX770,
     EX771,EX772,EX773,EX774,EX775,EX776,EX777,EX778,EX779,EX780,
     EX781,EX782,EX783,EX784,EX785,EX786,EX787,EX788,EX789,EX790,
     EX791,EX792,EX793,EX794,EX795,EX796,EX797,EX798,EX799,EX800,
     EX801,EX802,EX803,EX804,EX805,EX806,EX807,EX808,EX809,EX810,
     EX811,EX812,EX813,EX814,EX815,EX816,EX817,EX818,EX819,EX820,
     EX821,EX822,EX823,EX824,EX825,EX826,EX827,EX828,EX829,EX830,
     EX831,EX832,EX833,EX834,EX835,EX836,EX837,EX838,EX839,EX840,
     EX841,EX842,EX843,EX844,EX845,EX846,EX847,EX848,EX849,EX850,
     EX851,EX852,EX853,EX854,EX855,EX856,EX857,EX858,EX859,EX860,
     EX861,EX862,EX863,EX864,EX865,EX866,EX867,EX868,EX869,EX870,
     EX871,EX872,EX873,EX874,EX875,EX876,EX877,EX878,EX879,EX880,
     EX881,EX882,EX883,EX884,EX885,EX886,EX887,EX888,EX889,EX890,
     EX891,EX892,EX893,EX894,EX895,EX896,EX897,EX898,EX899,EX900,
     EX901,EX902,EX903,EX904,EX905,EX906,EX907,EX908,EX909,EX910,
     EX911,EX912,EX913,EX914,EX915,EX916,EX917,EX918,EX919,EX920,
     EX921,EX922,EX923,EX924,EX925,EX926,EX927,EX928,EX929,EX930,
     EX931,EX932,EX933,EX934,EX935,EX936,EX937,EX938,EX939,EX940,
     EX941,EX942,EX943,EX944,EX945,EX946,EX947,EX948,EX949,EX950,
     EX951,EX952,EX953,EX954,EX955,EX956,EX957,EX958,EX959,EX960,
     EX961,EX962,EX963,EX964,EX965,EX966,EX967,EX968,EX969,EX970,
     EX971,EX972,EX973,EX974,EX975,EX976,EX977,EX978,EX979,EX980,
     EX981,EX982,EX983,EX984,EX985,EX986,EX987,EX988,EX989,EX990,
     EX991,EX992,EX993,EX994,EX995,EX996,EX997,EX998,EX999,EX1000,
     EX1001,EX1002,EX1003,EX1004,EX1005,EX1006,EX1007,EX1008,EX1009,EX1010,
     EX1011,EX1012,EX1013,EX1014,EX1015,EX1016,EX1017,EX1018,EX1019,EX1020,
     EX1021,EX1022,EX1023,EX1024,EX1025,EX1026,EX1027,EX1028,EX1029,EX1030,
     EX1031,EX1032,EX1033,EX1034,EX1035,EX1036,EX1037,EX1038,EX1039,EX1040,
     EX1041,EX1042,EX1043,EX1044,EX1045,EX1046,EX1047,EX1048,EX1049,EX1050,
     EX1051,EX1052,EX1053,EX1054,EX1055,EX1056,EX1057,EX1058,EX1059,EX1060,
     EX1061,EX1062,EX1063,EX1064,EX1065,EX1066,EX1067,EX1068,EX1069,EX1070,
     EX1071,EX1072,EX1073,EX1074,EX1075,EX1076,EX1077,EX1078,EX1079,EX1080,
     EX1081,EX1082,EX1083,EX1084,EX1085,EX1086,EX1087,EX1088,EX1089,EX1090,
     EX1091,EX1092,EX1093,EX1094,EX1095,EX1096,EX1097,EX1098,EX1099,EX1100,
     EX1101,EX1102,EX1103,EX1104,EX1105,EX1106,EX1107,EX1108,EX1109,EX1110,
     EX1111,EX1112,EX1113,EX1114,EX1115,EX1116,EX1117,EX1118,EX1119,EX1120,
     EX1121,EX1122,EX1123,EX1124,EX1125,EX1126,EX1127,EX1128,EX1129,EX1130,
     EX1131,EX1132,EX1133,EX1134,EX1135,EX1136,EX1137,EX1138,EX1139,EX1140,
     EX1141,EX1142,EX1143,EX1144,EX1145,EX1146,EX1147,EX1148,EX1149,EX1150,
     EX1151,EX1152,EX1153,EX1154,EX1155,EX1156,EX1157,EX1158,EX1159,EX1160,
     EX1161,EX1162,EX1163,EX1164,EX1165,EX1166,EX1167,EX1168,EX1169,EX1170,
     EX1171,EX1172,EX1173,EX1174,EX1175,EX1176,EX1177,EX1178,EX1179,EX1180,
     EX1181,EX1182,EX1183,EX1184,EX1185,EX1186,EX1187,EX1188,EX1189,EX1190,
     EX1191,EX1192,EX1193,EX1194,EX1195,EX1196,EX1197,EX1198,EX1199,EX1200,
     EX1201,EX1202,EX1203,EX1204,EX1205,EX1206,EX1207,EX1208,EX1209,EX1210,
     EX1211,EX1212,EX1213,EX1214,EX1215,EX1216,EX1217,EX1218,EX1219,EX1220,
     EX1221,EX1222,EX1223,EX1224,EX1225,EX1226,EX1227,EX1228,EX1229,EX1230,
     EX1231,EX1232,EX1233,EX1234,EX1235,EX1236,EX1237,EX1238,EX1239,EX1240,
     EX1241,EX1242,EX1243,EX1244,EX1245,EX1246,EX1247,EX1248,EX1249,EX1250,
     EX1251,EX1252,EX1253,EX1254,EX1255,EX1256,EX1257,EX1258,EX1259,EX1260,
     EX1261,EX1262,EX1263,EX1264,EX1265,EX1266,EX1267,EX1268,EX1269,EX1270,
     EX1271,EX1272,EX1273,EX1274,EX1275,EX1276,EX1277,EX1278,EX1279,EX1280,
     EX1281,EX1282,EX1283,EX1284,EX1285,EX1286,EX1287,EX1288,EX1289,EX1290,
     EX1291,EX1292,EX1293,EX1294,EX1295,EX1296,EX1297,EX1298,EX1299,EX1300,
     EX1301,EX1302,EX1303,EX1304,EX1305,EX1306,EX1307,EX1308,EX1309,EX1310,
     EX1311,EX1312,EX1313,EX1314,EX1315,EX1316,EX1317,EX1318,EX1319,EX1320,
     EX1321,EX1322,EX1323,EX1324,EX1325,EX1326,EX1327,EX1328,EX1329,EX1330,
     EX1331,EX1332,EX1333,EX1334,EX1335,EX1336,EX1337,EX1338,EX1339,EX1340,
     EX1341,EX1342,EX1343,EX1344,EX1345,EX1346,EX1347,EX1348,EX1349,EX1350,
     EX1351,EX1352,EX1353,EX1354,EX1355,EX1356,EX1357,EX1358,EX1359,EX1360,
     EX1361,EX1362,EX1363,EX1364,EX1365,EX1366,EX1367,EX1368,EX1369,EX1370,
     EX1371,EX1372,EX1373,EX1374,EX1375,EX1376,EX1377,EX1378,EX1379,EX1380,
     EX1381,EX1382,EX1383,EX1384,EX1385,EX1386,EX1387,EX1388,EX1389,EX1390,
     EX1391,EX1392,EX1393,EX1394,EX1395,EX1396,EX1397,EX1398,EX1399,EX1400,
     EX1401,EX1402,EX1403,EX1404,EX1405,EX1406,EX1407,EX1408,EX1409,EX1410,
     EX1411,EX1412,EX1413,EX1414,EX1415,EX1416,EX1417,EX1418,EX1419,EX1420,
     EX1421,EX1422,EX1423,EX1424,EX1425,EX1426,EX1427,EX1428,EX1429,EX1430,
     EX1431,EX1432,EX1433,EX1434,EX1435,EX1436,EX1437,EX1438,EX1439,EX1440,
     EX1441,EX1442,EX1443,EX1444,EX1445,EX1446,EX1447,EX1448,EX1449,EX1450,
     EX1451,EX1452,EX1453,EX1454,EX1455,EX1456,EX1457,EX1458,EX1459,EX1460,
     EX1461,EX1462,EX1463,EX1464,EX1465,EX1466,EX1467,EX1468,EX1469,EX1470,
     EX1471,EX1472,EX1473,EX1474,EX1475,EX1476,EX1477,EX1478,EX1479,EX1480,
     EX1481,EX1482,EX1483,EX1484,EX1485,EX1486,EX1487,EX1488,EX1489,EX1490,
     EX1491,EX1492,EX1493,EX1494,EX1495,EX1496,EX1497,EX1498,EX1499,EX1500,
     EX1501,EX1502,EX1503,EX1504,EX1505,EX1506,EX1507,EX1508,EX1509,EX1510,
     EX1511,EX1512,EX1513,EX1514,EX1515,EX1516,EX1517,EX1518,EX1519,EX1520,
     EX1521,EX1522,EX1523,EX1524,EX1525,EX1526,EX1527,EX1528,EX1529,EX1530,
     EX1531,EX1532,EX1533,EX1534,EX1535,EX1536,EX1537,EX1538,EX1539,EX1540,
     EX1541,EX1542,EX1543,EX1544,EX1545,EX1546,EX1547,EX1548,EX1549,EX1550,
     EX1551,EX1552,EX1553,EX1554,EX1555,EX1556,EX1557,EX1558,EX1559,EX1560,
     EX1561,EX1562,EX1563,EX1564,EX1565,EX1566,EX1567,EX1568,EX1569,EX1570,
     EX1571,EX1572,EX1573,EX1574,EX1575,EX1576,EX1577,EX1578,EX1579,EX1580,
     EX1581,EX1582,EX1583,EX1584,EX1585,EX1586,EX1587,EX1588,EX1589,EX1590,
     EX1591,EX1592,EX1593,EX1594,EX1595,EX1596,EX1597,EX1598,EX1599,EX1600,
     EX1601,EX1602,EX1603,EX1604,EX1605,EX1606,EX1607,EX1608,EX1609,EX1610,
     EX1611,EX1612,EX1613,EX1614,EX1615,EX1616,EX1617,EX1618,EX1619,EX1620,
     EX1621,EX1622,EX1623,EX1624,EX1625,EX1626,EX1627,EX1628,EX1629,EX1630,
     EX1631,EX1632,EX1633,EX1634,EX1635,EX1636,EX1637,EX1638,EX1639,EX1640,N1,N13,N20,N33,N41,N45,N50,N58,N68,N77,N87,N97,N107,N116,N124,N125,N128,N132,N137,N143,N150,N159,N169,N179,N190,N200,N213,N222,N223,N226,N232,N238,N244,N250,N257,N264,N270,N274,N283,N294,N303,N311,N317,N322,N326,N329,N330,N343,N349,N350,N1713,N1947,N3195,N3833,N3987,N4028,N4145,N4589,N4667,N4815,N4944,N5002,N5045,N5047,N5078,N5102,N5120,N5121,N5192,N5231,N5360,N5361;


buf1 gate1( .a(N50), .O(N655) );
inv1 gate2( .a(N50), .O(N665) );
buf1 gate3( .a(N58), .O(N670) );
inv1 gate4( .a(N58), .O(N679) );
buf1 gate5( .a(N68), .O(N683) );
inv1 gate6( .a(N68), .O(N686) );
buf1 gate7( .a(N68), .O(N690) );
buf1 gate8( .a(N77), .O(N699) );
inv1 gate9( .a(N77), .O(N702) );
buf1 gate10( .a(N77), .O(N706) );
buf1 gate11( .a(N87), .O(N715) );
inv1 gate12( .a(N87), .O(N724) );
buf1 gate13( .a(N97), .O(N727) );
inv1 gate14( .a(N97), .O(N736) );
buf1 gate15( .a(N107), .O(N740) );
inv1 gate16( .a(N107), .O(N749) );
buf1 gate17( .a(N116), .O(N753) );
inv1 gate18( .a(N116), .O(N763) );
inv1 gate( .a(N257),.O(N257_NOT) );
inv1 gate( .a(N264),.O(N264_NOT));
and2 gate( .a(N257_NOT), .b(p1), .O(EX1) );
and2 gate( .a(N264_NOT), .b(EX1), .O(EX2) );
and2 gate( .a(N257), .b(p2), .O(EX3) );
and2 gate( .a(N264_NOT), .b(EX3), .O(EX4) );
and2 gate( .a(N257_NOT), .b(p3), .O(EX5) );
and2 gate( .a(N264), .b(EX5), .O(EX6) );
and2 gate( .a(N257), .b(p4), .O(EX7) );
and2 gate( .a(N264), .b(EX7), .O(EX8) );
or2  gate( .a(EX2), .b(EX4), .O(EX9) );
or2  gate( .a(EX6), .b(EX9), .O(EX10) );
or2  gate( .a(EX8), .b(EX10), .O(N768) );
inv1 gate20( .a(N1), .O(N769) );
buf1 gate21( .a(N1), .O(N772) );
inv1 gate22( .a(N1), .O(N779) );
buf1 gate23( .a(N13), .O(N782) );
inv1 gate24( .a(N13), .O(N786) );
inv1 gate( .a(N13),.O(N13_NOT) );
inv1 gate( .a(N20),.O(N20_NOT));
and2 gate( .a(N13_NOT), .b(p5), .O(EX11) );
and2 gate( .a(N20_NOT), .b(EX11), .O(EX12) );
and2 gate( .a(N13), .b(p6), .O(EX13) );
and2 gate( .a(N20_NOT), .b(EX13), .O(EX14) );
and2 gate( .a(N13_NOT), .b(p7), .O(EX15) );
and2 gate( .a(N20), .b(EX15), .O(EX16) );
and2 gate( .a(N13), .b(p8), .O(EX17) );
and2 gate( .a(N20), .b(EX17), .O(EX18) );
or2  gate( .a(EX12), .b(EX14), .O(EX19) );
or2  gate( .a(EX16), .b(EX19), .O(EX20) );
or2  gate( .a(EX18), .b(EX20), .O(N793) );
inv1 gate26( .a(N20), .O(N794) );
buf1 gate27( .a(N20), .O(N798) );
inv1 gate28( .a(N20), .O(N803) );
inv1 gate29( .a(N33), .O(N820) );
buf1 gate30( .a(N33), .O(N821) );
inv1 gate31( .a(N33), .O(N825) );
inv1 gate( .a(N33),.O(N33_NOT) );
inv1 gate( .a(N41),.O(N41_NOT));
and2 gate( .a(N33_NOT), .b(p9), .O(EX21) );
and2 gate( .a(N41_NOT), .b(EX21), .O(EX22) );
and2 gate( .a(N33), .b(p10), .O(EX23) );
and2 gate( .a(N41_NOT), .b(EX23), .O(EX24) );
and2 gate( .a(N33_NOT), .b(p11), .O(EX25) );
and2 gate( .a(N41), .b(EX25), .O(EX26) );
and2 gate( .a(N33), .b(p12), .O(EX27) );
and2 gate( .a(N41), .b(EX27), .O(EX28) );
or2  gate( .a(EX22), .b(EX24), .O(EX29) );
or2  gate( .a(EX26), .b(EX29), .O(EX30) );
or2  gate( .a(EX28), .b(EX30), .O(N829) );
inv1 gate33( .a(N41), .O(N832) );
inv1 gate( .a(N41),.O(N41_NOT) );
inv1 gate( .a(N45),.O(N45_NOT));
and2 gate( .a(N41_NOT), .b(p13), .O(EX31) );
and2 gate( .a(N45_NOT), .b(EX31), .O(EX32) );
and2 gate( .a(N41), .b(p14), .O(EX33) );
and2 gate( .a(N45_NOT), .b(EX33), .O(EX34) );
and2 gate( .a(N41_NOT), .b(p15), .O(EX35) );
and2 gate( .a(N45), .b(EX35), .O(EX36) );
and2 gate( .a(N41), .b(p16), .O(EX37) );
and2 gate( .a(N45), .b(EX37), .O(EX38) );
or2  gate( .a(EX32), .b(EX34), .O(EX39) );
or2  gate( .a(EX36), .b(EX39), .O(EX40) );
or2  gate( .a(EX38), .b(EX40), .O(N835) );
buf1 gate35( .a(N45), .O(N836) );
inv1 gate36( .a(N45), .O(N839) );
inv1 gate37( .a(N50), .O(N842) );
buf1 gate38( .a(N58), .O(N845) );
inv1 gate39( .a(N58), .O(N848) );
buf1 gate40( .a(N68), .O(N851) );
inv1 gate41( .a(N68), .O(N854) );
buf1 gate42( .a(N87), .O(N858) );
inv1 gate43( .a(N87), .O(N861) );
buf1 gate44( .a(N97), .O(N864) );
inv1 gate45( .a(N97), .O(N867) );
inv1 gate46( .a(N107), .O(N870) );
buf1 gate47( .a(N1), .O(N874) );
buf1 gate48( .a(N68), .O(N877) );
buf1 gate49( .a(N107), .O(N880) );
inv1 gate50( .a(N20), .O(N883) );
buf1 gate51( .a(N190), .O(N886) );
inv1 gate52( .a(N200), .O(N889) );
inv1 gate( .a(N20),.O(N20_NOT) );
inv1 gate( .a(N200),.O(N200_NOT));
and2 gate( .a(N20_NOT), .b(p17), .O(EX41) );
and2 gate( .a(N200_NOT), .b(EX41), .O(EX42) );
and2 gate( .a(N20), .b(p18), .O(EX43) );
and2 gate( .a(N200_NOT), .b(EX43), .O(EX44) );
and2 gate( .a(N20_NOT), .b(p19), .O(EX45) );
and2 gate( .a(N200), .b(EX45), .O(EX46) );
and2 gate( .a(N20), .b(p20), .O(EX47) );
and2 gate( .a(N200), .b(EX47), .O(EX48) );
or2  gate( .a(EX42), .b(EX44), .O(EX49) );
or2  gate( .a(EX46), .b(EX49), .O(EX50) );
or2  gate( .a(EX48), .b(EX50), .O(N890) );
inv1 gate( .a(N20),.O(N20_NOT) );
inv1 gate( .a(N200),.O(N200_NOT));
and2 gate( .a(N20_NOT), .b(p21), .O(EX51) );
and2 gate( .a(N200_NOT), .b(EX51), .O(EX52) );
and2 gate( .a(N20), .b(p22), .O(EX53) );
and2 gate( .a(N200_NOT), .b(EX53), .O(EX54) );
and2 gate( .a(N20_NOT), .b(p23), .O(EX55) );
and2 gate( .a(N200), .b(EX55), .O(EX56) );
and2 gate( .a(N20), .b(p24), .O(EX57) );
and2 gate( .a(N200), .b(EX57), .O(EX58) );
or2  gate( .a(EX52), .b(EX54), .O(EX59) );
or2  gate( .a(EX56), .b(EX59), .O(EX60) );
or2  gate( .a(EX58), .b(EX60), .O(N891) );
and2 gate55( .a(N20), .b(N179), .O(N892) );
inv1 gate56( .a(N20), .O(N895) );
inv1 gate( .a(N349),.O(N349_NOT) );
inv1 gate( .a(N33),.O(N33_NOT));
and2 gate( .a(N349_NOT), .b(p25), .O(EX61) );
and2 gate( .a(N33_NOT), .b(EX61), .O(EX62) );
and2 gate( .a(N349), .b(p26), .O(EX63) );
and2 gate( .a(N33_NOT), .b(EX63), .O(EX64) );
and2 gate( .a(N349_NOT), .b(p27), .O(EX65) );
and2 gate( .a(N33), .b(EX65), .O(EX66) );
and2 gate( .a(N349), .b(p28), .O(EX67) );
and2 gate( .a(N33), .b(EX67), .O(EX68) );
or2  gate( .a(EX62), .b(EX64), .O(EX69) );
or2  gate( .a(EX66), .b(EX69), .O(EX70) );
or2  gate( .a(EX68), .b(EX70), .O(N896) );
nand2 gate58( .a(N1), .b(N13), .O(N913) );
nand3 gate59( .a(N1), .b(N20), .c(N33), .O(N914) );
inv1 gate60( .a(N20), .O(N915) );
inv1 gate61( .a(N33), .O(N916) );
buf1 gate62( .a(N179), .O(N917) );
inv1 gate63( .a(N213), .O(N920) );
buf1 gate64( .a(N343), .O(N923) );
buf1 gate65( .a(N226), .O(N926) );
buf1 gate66( .a(N232), .O(N929) );
buf1 gate67( .a(N238), .O(N932) );
buf1 gate68( .a(N244), .O(N935) );
buf1 gate69( .a(N250), .O(N938) );
buf1 gate70( .a(N257), .O(N941) );
buf1 gate71( .a(N264), .O(N944) );
buf1 gate72( .a(N270), .O(N947) );
buf1 gate73( .a(N50), .O(N950) );
buf1 gate74( .a(N58), .O(N953) );
buf1 gate75( .a(N58), .O(N956) );
buf1 gate76( .a(N97), .O(N959) );
buf1 gate77( .a(N97), .O(N962) );
buf1 gate78( .a(N330), .O(N965) );
and2 gate79( .a(N250), .b(N768), .O(N1067) );
or2 gate80( .a(N820), .b(N20), .O(N1117) );
inv1 gate( .a(N895),.O(N895_NOT) );
inv1 gate( .a(N169),.O(N169_NOT));
and2 gate( .a(N895_NOT), .b(p29), .O(EX71) );
and2 gate( .a(N169_NOT), .b(EX71), .O(EX72) );
and2 gate( .a(N895), .b(p30), .O(EX73) );
and2 gate( .a(N169_NOT), .b(EX73), .O(EX74) );
and2 gate( .a(N895_NOT), .b(p31), .O(EX75) );
and2 gate( .a(N169), .b(EX75), .O(EX76) );
and2 gate( .a(N895), .b(p32), .O(EX77) );
and2 gate( .a(N169), .b(EX77), .O(EX78) );
or2  gate( .a(EX72), .b(EX74), .O(EX79) );
or2  gate( .a(EX76), .b(EX79), .O(EX80) );
or2  gate( .a(EX78), .b(EX80), .O(N1179) );
inv1 gate82( .a(N793), .O(N1196) );
inv1 gate( .a(N915),.O(N915_NOT) );
inv1 gate( .a(N1),.O(N1_NOT));
and2 gate( .a(N915_NOT), .b(p33), .O(EX81) );
and2 gate( .a(N1_NOT), .b(EX81), .O(EX82) );
and2 gate( .a(N915), .b(p34), .O(EX83) );
and2 gate( .a(N1_NOT), .b(EX83), .O(EX84) );
and2 gate( .a(N915_NOT), .b(p35), .O(EX85) );
and2 gate( .a(N1), .b(EX85), .O(EX86) );
and2 gate( .a(N915), .b(p36), .O(EX87) );
and2 gate( .a(N1), .b(EX87), .O(EX88) );
or2  gate( .a(EX82), .b(EX84), .O(EX89) );
or2  gate( .a(EX86), .b(EX89), .O(EX90) );
or2  gate( .a(EX88), .b(EX90), .O(N1197) );
and2 gate84( .a(N913), .b(N914), .O(N1202) );
inv1 gate( .a(N916),.O(N916_NOT) );
inv1 gate( .a(N1),.O(N1_NOT));
and2 gate( .a(N916_NOT), .b(p37), .O(EX91) );
and2 gate( .a(N1_NOT), .b(EX91), .O(EX92) );
and2 gate( .a(N916), .b(p38), .O(EX93) );
and2 gate( .a(N1_NOT), .b(EX93), .O(EX94) );
and2 gate( .a(N916_NOT), .b(p39), .O(EX95) );
and2 gate( .a(N1), .b(EX95), .O(EX96) );
and2 gate( .a(N916), .b(p40), .O(EX97) );
and2 gate( .a(N1), .b(EX97), .O(EX98) );
or2  gate( .a(EX92), .b(EX94), .O(EX99) );
or2  gate( .a(EX96), .b(EX99), .O(EX100) );
or2  gate( .a(EX98), .b(EX100), .O(N1219) );
and3 gate86( .a(N842), .b(N848), .c(N854), .O(N1250) );
inv1 gate( .a(N226),.O(N226_NOT) );
inv1 gate( .a(N655),.O(N655_NOT));
and2 gate( .a(N226_NOT), .b(p41), .O(EX101) );
and2 gate( .a(N655_NOT), .b(EX101), .O(EX102) );
and2 gate( .a(N226), .b(p42), .O(EX103) );
and2 gate( .a(N655_NOT), .b(EX103), .O(EX104) );
and2 gate( .a(N226_NOT), .b(p43), .O(EX105) );
and2 gate( .a(N655), .b(EX105), .O(EX106) );
and2 gate( .a(N226), .b(p44), .O(EX107) );
and2 gate( .a(N655), .b(EX107), .O(EX108) );
or2  gate( .a(EX102), .b(EX104), .O(EX109) );
or2  gate( .a(EX106), .b(EX109), .O(EX110) );
or2  gate( .a(EX108), .b(EX110), .O(N1251) );
inv1 gate( .a(N232),.O(N232_NOT) );
inv1 gate( .a(N670),.O(N670_NOT));
and2 gate( .a(N232_NOT), .b(p45), .O(EX111) );
and2 gate( .a(N670_NOT), .b(EX111), .O(EX112) );
and2 gate( .a(N232), .b(p46), .O(EX113) );
and2 gate( .a(N670_NOT), .b(EX113), .O(EX114) );
and2 gate( .a(N232_NOT), .b(p47), .O(EX115) );
and2 gate( .a(N670), .b(EX115), .O(EX116) );
and2 gate( .a(N232), .b(p48), .O(EX117) );
and2 gate( .a(N670), .b(EX117), .O(EX118) );
or2  gate( .a(EX112), .b(EX114), .O(EX119) );
or2  gate( .a(EX116), .b(EX119), .O(EX120) );
or2  gate( .a(EX118), .b(EX120), .O(N1252) );
nand2 gate89( .a(N238), .b(N690), .O(N1253) );
nand2 gate90( .a(N244), .b(N706), .O(N1254) );
inv1 gate( .a(N250),.O(N250_NOT) );
inv1 gate( .a(N715),.O(N715_NOT));
and2 gate( .a(N250_NOT), .b(p49), .O(EX121) );
and2 gate( .a(N715_NOT), .b(EX121), .O(EX122) );
and2 gate( .a(N250), .b(p50), .O(EX123) );
and2 gate( .a(N715_NOT), .b(EX123), .O(EX124) );
and2 gate( .a(N250_NOT), .b(p51), .O(EX125) );
and2 gate( .a(N715), .b(EX125), .O(EX126) );
and2 gate( .a(N250), .b(p52), .O(EX127) );
and2 gate( .a(N715), .b(EX127), .O(EX128) );
or2  gate( .a(EX122), .b(EX124), .O(EX129) );
or2  gate( .a(EX126), .b(EX129), .O(EX130) );
or2  gate( .a(EX128), .b(EX130), .O(N1255) );
inv1 gate( .a(N257),.O(N257_NOT) );
inv1 gate( .a(N727),.O(N727_NOT));
and2 gate( .a(N257_NOT), .b(p53), .O(EX131) );
and2 gate( .a(N727_NOT), .b(EX131), .O(EX132) );
and2 gate( .a(N257), .b(p54), .O(EX133) );
and2 gate( .a(N727_NOT), .b(EX133), .O(EX134) );
and2 gate( .a(N257_NOT), .b(p55), .O(EX135) );
and2 gate( .a(N727), .b(EX135), .O(EX136) );
and2 gate( .a(N257), .b(p56), .O(EX137) );
and2 gate( .a(N727), .b(EX137), .O(EX138) );
or2  gate( .a(EX132), .b(EX134), .O(EX139) );
or2  gate( .a(EX136), .b(EX139), .O(EX140) );
or2  gate( .a(EX138), .b(EX140), .O(N1256) );
inv1 gate( .a(N264),.O(N264_NOT) );
inv1 gate( .a(N740),.O(N740_NOT));
and2 gate( .a(N264_NOT), .b(p57), .O(EX141) );
and2 gate( .a(N740_NOT), .b(EX141), .O(EX142) );
and2 gate( .a(N264), .b(p58), .O(EX143) );
and2 gate( .a(N740_NOT), .b(EX143), .O(EX144) );
and2 gate( .a(N264_NOT), .b(p59), .O(EX145) );
and2 gate( .a(N740), .b(EX145), .O(EX146) );
and2 gate( .a(N264), .b(p60), .O(EX147) );
and2 gate( .a(N740), .b(EX147), .O(EX148) );
or2  gate( .a(EX142), .b(EX144), .O(EX149) );
or2  gate( .a(EX146), .b(EX149), .O(EX150) );
or2  gate( .a(EX148), .b(EX150), .O(N1257) );
nand2 gate94( .a(N270), .b(N753), .O(N1258) );
inv1 gate95( .a(N926), .O(N1259) );
inv1 gate96( .a(N929), .O(N1260) );
inv1 gate97( .a(N932), .O(N1261) );
inv1 gate98( .a(N935), .O(N1262) );
nand2 gate99( .a(N679), .b(N686), .O(N1263) );
nand2 gate100( .a(N736), .b(N749), .O(N1264) );
nand2 gate101( .a(N683), .b(N699), .O(N1267) );
buf1 gate102( .a(N665), .O(N1268) );
inv1 gate103( .a(N953), .O(N1271) );
inv1 gate104( .a(N959), .O(N1272) );
buf1 gate105( .a(N839), .O(N1273) );
buf1 gate106( .a(N839), .O(N1276) );
buf1 gate107( .a(N782), .O(N1279) );
buf1 gate108( .a(N825), .O(N1298) );
buf1 gate109( .a(N832), .O(N1302) );
and2 gate110( .a(N779), .b(N835), .O(N1306) );
and3 gate111( .a(N779), .b(N836), .c(N832), .O(N1315) );
and2 gate112( .a(N769), .b(N836), .O(N1322) );
and3 gate113( .a(N772), .b(N786), .c(N798), .O(N1325) );
nand3 gate114( .a(N772), .b(N786), .c(N798), .O(N1328) );
nand2 gate115( .a(N772), .b(N786), .O(N1331) );
buf1 gate116( .a(N874), .O(N1334) );
nand3 gate117( .a(N782), .b(N794), .c(N45), .O(N1337) );
nand3 gate118( .a(N842), .b(N848), .c(N854), .O(N1338) );
inv1 gate119( .a(N956), .O(N1339) );
and3 gate120( .a(N861), .b(N867), .c(N870), .O(N1340) );
nand3 gate121( .a(N861), .b(N867), .c(N870), .O(N1343) );
inv1 gate122( .a(N962), .O(N1344) );
inv1 gate123( .a(N803), .O(N1345) );
inv1 gate124( .a(N803), .O(N1346) );
inv1 gate125( .a(N803), .O(N1347) );
inv1 gate126( .a(N803), .O(N1348) );
inv1 gate127( .a(N803), .O(N1349) );
inv1 gate128( .a(N803), .O(N1350) );
inv1 gate129( .a(N803), .O(N1351) );
inv1 gate130( .a(N803), .O(N1352) );
or2 gate131( .a(N883), .b(N886), .O(N1353) );
nor2 gate132( .a(N883), .b(N886), .O(N1358) );
buf1 gate133( .a(N892), .O(N1363) );
inv1 gate134( .a(N892), .O(N1366) );
buf1 gate135( .a(N821), .O(N1369) );
buf1 gate136( .a(N825), .O(N1384) );
inv1 gate137( .a(N896), .O(N1401) );
inv1 gate138( .a(N896), .O(N1402) );
inv1 gate139( .a(N896), .O(N1403) );
inv1 gate140( .a(N896), .O(N1404) );
inv1 gate141( .a(N896), .O(N1405) );
inv1 gate142( .a(N896), .O(N1406) );
inv1 gate143( .a(N896), .O(N1407) );
inv1 gate144( .a(N896), .O(N1408) );
or2 gate145( .a(N1), .b(N1196), .O(N1409) );
inv1 gate146( .a(N829), .O(N1426) );
inv1 gate147( .a(N829), .O(N1427) );
and3 gate148( .a(N769), .b(N782), .c(N794), .O(N1452) );
inv1 gate149( .a(N917), .O(N1459) );
inv1 gate150( .a(N965), .O(N1460) );
inv1 gate( .a(N920),.O(N920_NOT) );
inv1 gate( .a(N923),.O(N923_NOT));
and2 gate( .a(N920_NOT), .b(p61), .O(EX151) );
and2 gate( .a(N923_NOT), .b(EX151), .O(EX152) );
and2 gate( .a(N920), .b(p62), .O(EX153) );
and2 gate( .a(N923_NOT), .b(EX153), .O(EX154) );
and2 gate( .a(N920_NOT), .b(p63), .O(EX155) );
and2 gate( .a(N923), .b(EX155), .O(EX156) );
and2 gate( .a(N920), .b(p64), .O(EX157) );
and2 gate( .a(N923), .b(EX157), .O(EX158) );
or2  gate( .a(EX152), .b(EX154), .O(EX159) );
or2  gate( .a(EX156), .b(EX159), .O(EX160) );
or2  gate( .a(EX158), .b(EX160), .O(N1461) );
inv1 gate( .a(N920),.O(N920_NOT) );
inv1 gate( .a(N923),.O(N923_NOT));
and2 gate( .a(N920_NOT), .b(p65), .O(EX161) );
and2 gate( .a(N923_NOT), .b(EX161), .O(EX162) );
and2 gate( .a(N920), .b(p66), .O(EX163) );
and2 gate( .a(N923_NOT), .b(EX163), .O(EX164) );
and2 gate( .a(N920_NOT), .b(p67), .O(EX165) );
and2 gate( .a(N923), .b(EX165), .O(EX166) );
and2 gate( .a(N920), .b(p68), .O(EX167) );
and2 gate( .a(N923), .b(EX167), .O(EX168) );
or2  gate( .a(EX162), .b(EX164), .O(EX169) );
or2  gate( .a(EX166), .b(EX169), .O(EX170) );
or2  gate( .a(EX168), .b(EX170), .O(N1464) );
inv1 gate153( .a(N938), .O(N1467) );
inv1 gate154( .a(N941), .O(N1468) );
inv1 gate155( .a(N944), .O(N1469) );
inv1 gate156( .a(N947), .O(N1470) );
buf1 gate157( .a(N679), .O(N1471) );
inv1 gate158( .a(N950), .O(N1474) );
buf1 gate159( .a(N686), .O(N1475) );
buf1 gate160( .a(N702), .O(N1478) );
buf1 gate161( .a(N724), .O(N1481) );
buf1 gate162( .a(N736), .O(N1484) );
buf1 gate163( .a(N749), .O(N1487) );
buf1 gate164( .a(N763), .O(N1490) );
buf1 gate165( .a(N877), .O(N1493) );
buf1 gate166( .a(N877), .O(N1496) );
buf1 gate167( .a(N880), .O(N1499) );
buf1 gate168( .a(N880), .O(N1502) );
inv1 gate( .a(N702),.O(N702_NOT) );
inv1 gate( .a(N1250),.O(N1250_NOT));
and2 gate( .a(N702_NOT), .b(p69), .O(EX171) );
and2 gate( .a(N1250_NOT), .b(EX171), .O(EX172) );
and2 gate( .a(N702), .b(p70), .O(EX173) );
and2 gate( .a(N1250_NOT), .b(EX173), .O(EX174) );
and2 gate( .a(N702_NOT), .b(p71), .O(EX175) );
and2 gate( .a(N1250), .b(EX175), .O(EX176) );
and2 gate( .a(N702), .b(p72), .O(EX177) );
and2 gate( .a(N1250), .b(EX177), .O(EX178) );
or2  gate( .a(EX172), .b(EX174), .O(EX179) );
or2  gate( .a(EX176), .b(EX179), .O(EX180) );
or2  gate( .a(EX178), .b(EX180), .O(N1505) );
and4 gate170( .a(N1251), .b(N1252), .c(N1253), .d(N1254), .O(N1507) );
and4 gate171( .a(N1255), .b(N1256), .c(N1257), .d(N1258), .O(N1508) );
nand2 gate172( .a(N929), .b(N1259), .O(N1509) );
nand2 gate173( .a(N926), .b(N1260), .O(N1510) );
nand2 gate174( .a(N935), .b(N1261), .O(N1511) );
nand2 gate175( .a(N932), .b(N1262), .O(N1512) );
and2 gate176( .a(N655), .b(N1263), .O(N1520) );
and2 gate177( .a(N874), .b(N1337), .O(N1562) );
inv1 gate178( .a(N1117), .O(N1579) );
and2 gate179( .a(N803), .b(N1117), .O(N1580) );
and2 gate180( .a(N1338), .b(N1345), .O(N1581) );
inv1 gate181( .a(N1117), .O(N1582) );
and2 gate182( .a(N803), .b(N1117), .O(N1583) );
inv1 gate183( .a(N1117), .O(N1584) );
and2 gate184( .a(N803), .b(N1117), .O(N1585) );
and2 gate185( .a(N854), .b(N1347), .O(N1586) );
inv1 gate186( .a(N1117), .O(N1587) );
and2 gate187( .a(N803), .b(N1117), .O(N1588) );
inv1 gate( .a(N77),.O(N77_NOT) );
inv1 gate( .a(N1348),.O(N1348_NOT));
and2 gate( .a(N77_NOT), .b(p73), .O(EX181) );
and2 gate( .a(N1348_NOT), .b(EX181), .O(EX182) );
and2 gate( .a(N77), .b(p74), .O(EX183) );
and2 gate( .a(N1348_NOT), .b(EX183), .O(EX184) );
and2 gate( .a(N77_NOT), .b(p75), .O(EX185) );
and2 gate( .a(N1348), .b(EX185), .O(EX186) );
and2 gate( .a(N77), .b(p76), .O(EX187) );
and2 gate( .a(N1348), .b(EX187), .O(EX188) );
or2  gate( .a(EX182), .b(EX184), .O(EX189) );
or2  gate( .a(EX186), .b(EX189), .O(EX190) );
or2  gate( .a(EX188), .b(EX190), .O(N1589) );
inv1 gate189( .a(N1117), .O(N1590) );
and2 gate190( .a(N803), .b(N1117), .O(N1591) );
and2 gate191( .a(N1343), .b(N1349), .O(N1592) );
inv1 gate192( .a(N1117), .O(N1593) );
inv1 gate( .a(N803),.O(N803_NOT) );
inv1 gate( .a(N1117),.O(N1117_NOT));
and2 gate( .a(N803_NOT), .b(p77), .O(EX191) );
and2 gate( .a(N1117_NOT), .b(EX191), .O(EX192) );
and2 gate( .a(N803), .b(p78), .O(EX193) );
and2 gate( .a(N1117_NOT), .b(EX193), .O(EX194) );
and2 gate( .a(N803_NOT), .b(p79), .O(EX195) );
and2 gate( .a(N1117), .b(EX195), .O(EX196) );
and2 gate( .a(N803), .b(p80), .O(EX197) );
and2 gate( .a(N1117), .b(EX197), .O(EX198) );
or2  gate( .a(EX192), .b(EX194), .O(EX199) );
or2  gate( .a(EX196), .b(EX199), .O(EX200) );
or2  gate( .a(EX198), .b(EX200), .O(N1594) );
inv1 gate194( .a(N1117), .O(N1595) );
and2 gate195( .a(N803), .b(N1117), .O(N1596) );
and2 gate196( .a(N870), .b(N1351), .O(N1597) );
inv1 gate197( .a(N1117), .O(N1598) );
and2 gate198( .a(N803), .b(N1117), .O(N1599) );
and2 gate199( .a(N116), .b(N1352), .O(N1600) );
and2 gate200( .a(N222), .b(N1401), .O(N1643) );
and2 gate201( .a(N223), .b(N1402), .O(N1644) );
and2 gate202( .a(N226), .b(N1403), .O(N1645) );
and2 gate203( .a(N232), .b(N1404), .O(N1646) );
inv1 gate( .a(N238),.O(N238_NOT) );
inv1 gate( .a(N1405),.O(N1405_NOT));
and2 gate( .a(N238_NOT), .b(p81), .O(EX201) );
and2 gate( .a(N1405_NOT), .b(EX201), .O(EX202) );
and2 gate( .a(N238), .b(p82), .O(EX203) );
and2 gate( .a(N1405_NOT), .b(EX203), .O(EX204) );
and2 gate( .a(N238_NOT), .b(p83), .O(EX205) );
and2 gate( .a(N1405), .b(EX205), .O(EX206) );
and2 gate( .a(N238), .b(p84), .O(EX207) );
and2 gate( .a(N1405), .b(EX207), .O(EX208) );
or2  gate( .a(EX202), .b(EX204), .O(EX209) );
or2  gate( .a(EX206), .b(EX209), .O(EX210) );
or2  gate( .a(EX208), .b(EX210), .O(N1647) );
inv1 gate( .a(N244),.O(N244_NOT) );
inv1 gate( .a(N1406),.O(N1406_NOT));
and2 gate( .a(N244_NOT), .b(p85), .O(EX211) );
and2 gate( .a(N1406_NOT), .b(EX211), .O(EX212) );
and2 gate( .a(N244), .b(p86), .O(EX213) );
and2 gate( .a(N1406_NOT), .b(EX213), .O(EX214) );
and2 gate( .a(N244_NOT), .b(p87), .O(EX215) );
and2 gate( .a(N1406), .b(EX215), .O(EX216) );
and2 gate( .a(N244), .b(p88), .O(EX217) );
and2 gate( .a(N1406), .b(EX217), .O(EX218) );
or2  gate( .a(EX212), .b(EX214), .O(EX219) );
or2  gate( .a(EX216), .b(EX219), .O(EX220) );
or2  gate( .a(EX218), .b(EX220), .O(N1648) );
and2 gate206( .a(N250), .b(N1407), .O(N1649) );
inv1 gate( .a(N257),.O(N257_NOT) );
inv1 gate( .a(N1408),.O(N1408_NOT));
and2 gate( .a(N257_NOT), .b(p89), .O(EX221) );
and2 gate( .a(N1408_NOT), .b(EX221), .O(EX222) );
and2 gate( .a(N257), .b(p90), .O(EX223) );
and2 gate( .a(N1408_NOT), .b(EX223), .O(EX224) );
and2 gate( .a(N257_NOT), .b(p91), .O(EX225) );
and2 gate( .a(N1408), .b(EX225), .O(EX226) );
and2 gate( .a(N257), .b(p92), .O(EX227) );
and2 gate( .a(N1408), .b(EX227), .O(EX228) );
or2  gate( .a(EX222), .b(EX224), .O(EX229) );
or2  gate( .a(EX226), .b(EX229), .O(EX230) );
or2  gate( .a(EX228), .b(EX230), .O(N1650) );
and3 gate208( .a(N1), .b(N13), .c(N1426), .O(N1667) );
and3 gate209( .a(N1), .b(N13), .c(N1427), .O(N1670) );
inv1 gate210( .a(N1202), .O(N1673) );
inv1 gate211( .a(N1202), .O(N1674) );
inv1 gate212( .a(N1202), .O(N1675) );
inv1 gate213( .a(N1202), .O(N1676) );
inv1 gate214( .a(N1202), .O(N1677) );
inv1 gate215( .a(N1202), .O(N1678) );
inv1 gate216( .a(N1202), .O(N1679) );
inv1 gate217( .a(N1202), .O(N1680) );
nand2 gate218( .a(N941), .b(N1467), .O(N1691) );
nand2 gate219( .a(N938), .b(N1468), .O(N1692) );
nand2 gate220( .a(N947), .b(N1469), .O(N1693) );
nand2 gate221( .a(N944), .b(N1470), .O(N1694) );
inv1 gate222( .a(N1505), .O(N1713) );
and2 gate223( .a(N87), .b(N1264), .O(N1714) );
nand2 gate224( .a(N1509), .b(N1510), .O(N1715) );
nand2 gate225( .a(N1511), .b(N1512), .O(N1718) );
nand2 gate226( .a(N1507), .b(N1508), .O(N1721) );
and2 gate227( .a(N763), .b(N1340), .O(N1722) );
nand2 gate228( .a(N763), .b(N1340), .O(N1725) );
inv1 gate229( .a(N1268), .O(N1726) );
nand2 gate230( .a(N1493), .b(N1271), .O(N1727) );
inv1 gate231( .a(N1493), .O(N1728) );
and2 gate232( .a(N683), .b(N1268), .O(N1729) );
nand2 gate233( .a(N1499), .b(N1272), .O(N1730) );
inv1 gate234( .a(N1499), .O(N1731) );
nand2 gate235( .a(N87), .b(N1264), .O(N1735) );
inv1 gate236( .a(N1273), .O(N1736) );
inv1 gate237( .a(N1276), .O(N1737) );
nand2 gate238( .a(N1325), .b(N821), .O(N1738) );
nand2 gate239( .a(N1325), .b(N825), .O(N1747) );
nand3 gate240( .a(N772), .b(N1279), .c(N798), .O(N1756) );
nand4 gate241( .a(N772), .b(N786), .c(N798), .d(N1302), .O(N1761) );
nand2 gate242( .a(N1496), .b(N1339), .O(N1764) );
inv1 gate243( .a(N1496), .O(N1765) );
inv1 gate( .a(N1502),.O(N1502_NOT) );
inv1 gate( .a(N1344),.O(N1344_NOT));
and2 gate( .a(N1502_NOT), .b(p93), .O(EX231) );
and2 gate( .a(N1344_NOT), .b(EX231), .O(EX232) );
and2 gate( .a(N1502), .b(p94), .O(EX233) );
and2 gate( .a(N1344_NOT), .b(EX233), .O(EX234) );
and2 gate( .a(N1502_NOT), .b(p95), .O(EX235) );
and2 gate( .a(N1344), .b(EX235), .O(EX236) );
and2 gate( .a(N1502), .b(p96), .O(EX237) );
and2 gate( .a(N1344), .b(EX237), .O(EX238) );
or2  gate( .a(EX232), .b(EX234), .O(EX239) );
or2  gate( .a(EX236), .b(EX239), .O(EX240) );
or2  gate( .a(EX238), .b(EX240), .O(N1766) );
inv1 gate245( .a(N1502), .O(N1767) );
inv1 gate246( .a(N1328), .O(N1768) );
inv1 gate247( .a(N1334), .O(N1769) );
inv1 gate248( .a(N1331), .O(N1770) );
and2 gate249( .a(N845), .b(N1579), .O(N1787) );
inv1 gate( .a(N150),.O(N150_NOT) );
inv1 gate( .a(N1580),.O(N1580_NOT));
and2 gate( .a(N150_NOT), .b(p97), .O(EX241) );
and2 gate( .a(N1580_NOT), .b(EX241), .O(EX242) );
and2 gate( .a(N150), .b(p98), .O(EX243) );
and2 gate( .a(N1580_NOT), .b(EX243), .O(EX244) );
and2 gate( .a(N150_NOT), .b(p99), .O(EX245) );
and2 gate( .a(N1580), .b(EX245), .O(EX246) );
and2 gate( .a(N150), .b(p100), .O(EX247) );
and2 gate( .a(N1580), .b(EX247), .O(EX248) );
or2  gate( .a(EX242), .b(EX244), .O(EX249) );
or2  gate( .a(EX246), .b(EX249), .O(EX250) );
or2  gate( .a(EX248), .b(EX250), .O(N1788) );
inv1 gate( .a(N851),.O(N851_NOT) );
inv1 gate( .a(N1582),.O(N1582_NOT));
and2 gate( .a(N851_NOT), .b(p101), .O(EX251) );
and2 gate( .a(N1582_NOT), .b(EX251), .O(EX252) );
and2 gate( .a(N851), .b(p102), .O(EX253) );
and2 gate( .a(N1582_NOT), .b(EX253), .O(EX254) );
and2 gate( .a(N851_NOT), .b(p103), .O(EX255) );
and2 gate( .a(N1582), .b(EX255), .O(EX256) );
and2 gate( .a(N851), .b(p104), .O(EX257) );
and2 gate( .a(N1582), .b(EX257), .O(EX258) );
or2  gate( .a(EX252), .b(EX254), .O(EX259) );
or2  gate( .a(EX256), .b(EX259), .O(EX260) );
or2  gate( .a(EX258), .b(EX260), .O(N1789) );
and2 gate252( .a(N159), .b(N1583), .O(N1790) );
and2 gate253( .a(N77), .b(N1584), .O(N1791) );
and2 gate254( .a(N50), .b(N1585), .O(N1792) );
inv1 gate( .a(N858),.O(N858_NOT) );
inv1 gate( .a(N1587),.O(N1587_NOT));
and2 gate( .a(N858_NOT), .b(p105), .O(EX261) );
and2 gate( .a(N1587_NOT), .b(EX261), .O(EX262) );
and2 gate( .a(N858), .b(p106), .O(EX263) );
and2 gate( .a(N1587_NOT), .b(EX263), .O(EX264) );
and2 gate( .a(N858_NOT), .b(p107), .O(EX265) );
and2 gate( .a(N1587), .b(EX265), .O(EX266) );
and2 gate( .a(N858), .b(p108), .O(EX267) );
and2 gate( .a(N1587), .b(EX267), .O(EX268) );
or2  gate( .a(EX262), .b(EX264), .O(EX269) );
or2  gate( .a(EX266), .b(EX269), .O(EX270) );
or2  gate( .a(EX268), .b(EX270), .O(N1793) );
and2 gate256( .a(N845), .b(N1588), .O(N1794) );
and2 gate257( .a(N864), .b(N1590), .O(N1795) );
and2 gate258( .a(N851), .b(N1591), .O(N1796) );
and2 gate259( .a(N107), .b(N1593), .O(N1797) );
and2 gate260( .a(N77), .b(N1594), .O(N1798) );
and2 gate261( .a(N116), .b(N1595), .O(N1799) );
and2 gate262( .a(N858), .b(N1596), .O(N1800) );
and2 gate263( .a(N283), .b(N1598), .O(N1801) );
and2 gate264( .a(N864), .b(N1599), .O(N1802) );
and2 gate265( .a(N200), .b(N1363), .O(N1803) );
and2 gate266( .a(N889), .b(N1363), .O(N1806) );
and2 gate267( .a(N890), .b(N1366), .O(N1809) );
inv1 gate( .a(N891),.O(N891_NOT) );
inv1 gate( .a(N1366),.O(N1366_NOT));
and2 gate( .a(N891_NOT), .b(p109), .O(EX271) );
and2 gate( .a(N1366_NOT), .b(EX271), .O(EX272) );
and2 gate( .a(N891), .b(p110), .O(EX273) );
and2 gate( .a(N1366_NOT), .b(EX273), .O(EX274) );
and2 gate( .a(N891_NOT), .b(p111), .O(EX275) );
and2 gate( .a(N1366), .b(EX275), .O(EX276) );
and2 gate( .a(N891), .b(p112), .O(EX277) );
and2 gate( .a(N1366), .b(EX277), .O(EX278) );
or2  gate( .a(EX272), .b(EX274), .O(EX279) );
or2  gate( .a(EX276), .b(EX279), .O(EX280) );
or2  gate( .a(EX278), .b(EX280), .O(N1812) );
nand2 gate269( .a(N1298), .b(N1302), .O(N1815) );
nand2 gate270( .a(N821), .b(N1302), .O(N1818) );
nand3 gate271( .a(N772), .b(N1279), .c(N1179), .O(N1821) );
nand3 gate272( .a(N786), .b(N794), .c(N1298), .O(N1824) );
inv1 gate( .a(N786),.O(N786_NOT) );
inv1 gate( .a(N1298),.O(N1298_NOT));
and2 gate( .a(N786_NOT), .b(p113), .O(EX281) );
and2 gate( .a(N1298_NOT), .b(EX281), .O(EX282) );
and2 gate( .a(N786), .b(p114), .O(EX283) );
and2 gate( .a(N1298_NOT), .b(EX283), .O(EX284) );
and2 gate( .a(N786_NOT), .b(p115), .O(EX285) );
and2 gate( .a(N1298), .b(EX285), .O(EX286) );
and2 gate( .a(N786), .b(p116), .O(EX287) );
and2 gate( .a(N1298), .b(EX287), .O(EX288) );
or2  gate( .a(EX282), .b(EX284), .O(EX289) );
or2  gate( .a(EX286), .b(EX289), .O(EX290) );
or2  gate( .a(EX288), .b(EX290), .O(N1833) );
inv1 gate274( .a(N1369), .O(N1842) );
inv1 gate275( .a(N1369), .O(N1843) );
inv1 gate276( .a(N1369), .O(N1844) );
inv1 gate277( .a(N1369), .O(N1845) );
inv1 gate278( .a(N1369), .O(N1846) );
inv1 gate279( .a(N1369), .O(N1847) );
inv1 gate280( .a(N1369), .O(N1848) );
inv1 gate281( .a(N1384), .O(N1849) );
and2 gate282( .a(N1384), .b(N896), .O(N1850) );
inv1 gate283( .a(N1384), .O(N1851) );
and2 gate284( .a(N1384), .b(N896), .O(N1852) );
inv1 gate285( .a(N1384), .O(N1853) );
and2 gate286( .a(N1384), .b(N896), .O(N1854) );
inv1 gate287( .a(N1384), .O(N1855) );
and2 gate288( .a(N1384), .b(N896), .O(N1856) );
inv1 gate289( .a(N1384), .O(N1857) );
and2 gate290( .a(N1384), .b(N896), .O(N1858) );
inv1 gate291( .a(N1384), .O(N1859) );
and2 gate292( .a(N1384), .b(N896), .O(N1860) );
inv1 gate293( .a(N1384), .O(N1861) );
and2 gate294( .a(N1384), .b(N896), .O(N1862) );
inv1 gate295( .a(N1384), .O(N1863) );
and2 gate296( .a(N1384), .b(N896), .O(N1864) );
and2 gate297( .a(N1202), .b(N1409), .O(N1869) );
nor2 gate298( .a(N50), .b(N1409), .O(N1870) );
inv1 gate299( .a(N1306), .O(N1873) );
and2 gate300( .a(N1202), .b(N1409), .O(N1874) );
nor2 gate301( .a(N58), .b(N1409), .O(N1875) );
inv1 gate302( .a(N1306), .O(N1878) );
and2 gate303( .a(N1202), .b(N1409), .O(N1879) );
inv1 gate( .a(N68),.O(N68_NOT) );
inv1 gate( .a(N1409),.O(N1409_NOT));
and2 gate( .a(N68_NOT), .b(p117), .O(EX291) );
and2 gate( .a(N1409_NOT), .b(EX291), .O(EX292) );
and2 gate( .a(N68), .b(p118), .O(EX293) );
and2 gate( .a(N1409_NOT), .b(EX293), .O(EX294) );
and2 gate( .a(N68_NOT), .b(p119), .O(EX295) );
and2 gate( .a(N1409), .b(EX295), .O(EX296) );
and2 gate( .a(N68), .b(p120), .O(EX297) );
and2 gate( .a(N1409), .b(EX297), .O(EX298) );
or2  gate( .a(EX292), .b(EX294), .O(EX299) );
or2  gate( .a(EX296), .b(EX299), .O(EX300) );
or2  gate( .a(EX298), .b(EX300), .O(N1880) );
inv1 gate305( .a(N1306), .O(N1883) );
and2 gate306( .a(N1202), .b(N1409), .O(N1884) );
nor2 gate307( .a(N77), .b(N1409), .O(N1885) );
inv1 gate308( .a(N1306), .O(N1888) );
and2 gate309( .a(N1202), .b(N1409), .O(N1889) );
nor2 gate310( .a(N87), .b(N1409), .O(N1890) );
inv1 gate311( .a(N1322), .O(N1893) );
inv1 gate( .a(N1202),.O(N1202_NOT) );
inv1 gate( .a(N1409),.O(N1409_NOT));
and2 gate( .a(N1202_NOT), .b(p121), .O(EX301) );
and2 gate( .a(N1409_NOT), .b(EX301), .O(EX302) );
and2 gate( .a(N1202), .b(p122), .O(EX303) );
and2 gate( .a(N1409_NOT), .b(EX303), .O(EX304) );
and2 gate( .a(N1202_NOT), .b(p123), .O(EX305) );
and2 gate( .a(N1409), .b(EX305), .O(EX306) );
and2 gate( .a(N1202), .b(p124), .O(EX307) );
and2 gate( .a(N1409), .b(EX307), .O(EX308) );
or2  gate( .a(EX302), .b(EX304), .O(EX309) );
or2  gate( .a(EX306), .b(EX309), .O(EX310) );
or2  gate( .a(EX308), .b(EX310), .O(N1894) );
nor2 gate313( .a(N97), .b(N1409), .O(N1895) );
inv1 gate314( .a(N1315), .O(N1898) );
inv1 gate( .a(N1202),.O(N1202_NOT) );
inv1 gate( .a(N1409),.O(N1409_NOT));
and2 gate( .a(N1202_NOT), .b(p125), .O(EX311) );
and2 gate( .a(N1409_NOT), .b(EX311), .O(EX312) );
and2 gate( .a(N1202), .b(p126), .O(EX313) );
and2 gate( .a(N1409_NOT), .b(EX313), .O(EX314) );
and2 gate( .a(N1202_NOT), .b(p127), .O(EX315) );
and2 gate( .a(N1409), .b(EX315), .O(EX316) );
and2 gate( .a(N1202), .b(p128), .O(EX317) );
and2 gate( .a(N1409), .b(EX317), .O(EX318) );
or2  gate( .a(EX312), .b(EX314), .O(EX319) );
or2  gate( .a(EX316), .b(EX319), .O(EX320) );
or2  gate( .a(EX318), .b(EX320), .O(N1899) );
nor2 gate316( .a(N107), .b(N1409), .O(N1900) );
inv1 gate317( .a(N1315), .O(N1903) );
and2 gate318( .a(N1202), .b(N1409), .O(N1904) );
nor2 gate319( .a(N116), .b(N1409), .O(N1905) );
inv1 gate320( .a(N1315), .O(N1908) );
and2 gate321( .a(N1452), .b(N213), .O(N1909) );
nand2 gate322( .a(N1452), .b(N213), .O(N1912) );
and3 gate323( .a(N1452), .b(N213), .c(N343), .O(N1913) );
nand3 gate324( .a(N1452), .b(N213), .c(N343), .O(N1917) );
and3 gate325( .a(N1452), .b(N213), .c(N343), .O(N1922) );
nand3 gate326( .a(N1452), .b(N213), .c(N343), .O(N1926) );
buf1 gate327( .a(N1464), .O(N1930) );
nand2 gate328( .a(N1691), .b(N1692), .O(N1933) );
inv1 gate( .a(N1693),.O(N1693_NOT) );
inv1 gate( .a(N1694),.O(N1694_NOT));
and2 gate( .a(N1693_NOT), .b(p129), .O(EX321) );
and2 gate( .a(N1694_NOT), .b(EX321), .O(EX322) );
and2 gate( .a(N1693), .b(p130), .O(EX323) );
and2 gate( .a(N1694_NOT), .b(EX323), .O(EX324) );
and2 gate( .a(N1693_NOT), .b(p131), .O(EX325) );
and2 gate( .a(N1694), .b(EX325), .O(EX326) );
and2 gate( .a(N1693), .b(p132), .O(EX327) );
and2 gate( .a(N1694), .b(EX327), .O(EX328) );
or2  gate( .a(EX322), .b(EX324), .O(EX329) );
or2  gate( .a(EX326), .b(EX329), .O(EX330) );
or2  gate( .a(EX328), .b(EX330), .O(N1936) );
inv1 gate330( .a(N1471), .O(N1939) );
nand2 gate331( .a(N1471), .b(N1474), .O(N1940) );
inv1 gate332( .a(N1475), .O(N1941) );
inv1 gate333( .a(N1478), .O(N1942) );
inv1 gate334( .a(N1481), .O(N1943) );
inv1 gate335( .a(N1484), .O(N1944) );
inv1 gate336( .a(N1487), .O(N1945) );
inv1 gate337( .a(N1490), .O(N1946) );
inv1 gate338( .a(N1714), .O(N1947) );
nand2 gate339( .a(N953), .b(N1728), .O(N1960) );
nand2 gate340( .a(N959), .b(N1731), .O(N1961) );
and2 gate341( .a(N1520), .b(N1276), .O(N1966) );
nand2 gate342( .a(N956), .b(N1765), .O(N1981) );
nand2 gate343( .a(N962), .b(N1767), .O(N1982) );
and2 gate344( .a(N1067), .b(N1768), .O(N1983) );
or3 gate345( .a(N1581), .b(N1787), .c(N1788), .O(N1986) );
or3 gate346( .a(N1586), .b(N1791), .c(N1792), .O(N1987) );
or3 gate347( .a(N1589), .b(N1793), .c(N1794), .O(N1988) );
or3 gate348( .a(N1592), .b(N1795), .c(N1796), .O(N1989) );
or3 gate349( .a(N1597), .b(N1799), .c(N1800), .O(N1990) );
or3 gate350( .a(N1600), .b(N1801), .c(N1802), .O(N1991) );
and2 gate351( .a(N77), .b(N1849), .O(N2022) );
inv1 gate( .a(N223),.O(N223_NOT) );
inv1 gate( .a(N1850),.O(N1850_NOT));
and2 gate( .a(N223_NOT), .b(p133), .O(EX331) );
and2 gate( .a(N1850_NOT), .b(EX331), .O(EX332) );
and2 gate( .a(N223), .b(p134), .O(EX333) );
and2 gate( .a(N1850_NOT), .b(EX333), .O(EX334) );
and2 gate( .a(N223_NOT), .b(p135), .O(EX335) );
and2 gate( .a(N1850), .b(EX335), .O(EX336) );
and2 gate( .a(N223), .b(p136), .O(EX337) );
and2 gate( .a(N1850), .b(EX337), .O(EX338) );
or2  gate( .a(EX332), .b(EX334), .O(EX339) );
or2  gate( .a(EX336), .b(EX339), .O(EX340) );
or2  gate( .a(EX338), .b(EX340), .O(N2023) );
and2 gate353( .a(N87), .b(N1851), .O(N2024) );
and2 gate354( .a(N226), .b(N1852), .O(N2025) );
and2 gate355( .a(N97), .b(N1853), .O(N2026) );
and2 gate356( .a(N232), .b(N1854), .O(N2027) );
inv1 gate( .a(N107),.O(N107_NOT) );
inv1 gate( .a(N1855),.O(N1855_NOT));
and2 gate( .a(N107_NOT), .b(p137), .O(EX341) );
and2 gate( .a(N1855_NOT), .b(EX341), .O(EX342) );
and2 gate( .a(N107), .b(p138), .O(EX343) );
and2 gate( .a(N1855_NOT), .b(EX343), .O(EX344) );
and2 gate( .a(N107_NOT), .b(p139), .O(EX345) );
and2 gate( .a(N1855), .b(EX345), .O(EX346) );
and2 gate( .a(N107), .b(p140), .O(EX347) );
and2 gate( .a(N1855), .b(EX347), .O(EX348) );
or2  gate( .a(EX342), .b(EX344), .O(EX349) );
or2  gate( .a(EX346), .b(EX349), .O(EX350) );
or2  gate( .a(EX348), .b(EX350), .O(N2028) );
and2 gate358( .a(N238), .b(N1856), .O(N2029) );
and2 gate359( .a(N116), .b(N1857), .O(N2030) );
and2 gate360( .a(N244), .b(N1858), .O(N2031) );
and2 gate361( .a(N283), .b(N1859), .O(N2032) );
and2 gate362( .a(N250), .b(N1860), .O(N2033) );
and2 gate363( .a(N294), .b(N1861), .O(N2034) );
and2 gate364( .a(N257), .b(N1862), .O(N2035) );
inv1 gate( .a(N303),.O(N303_NOT) );
inv1 gate( .a(N1863),.O(N1863_NOT));
and2 gate( .a(N303_NOT), .b(p141), .O(EX351) );
and2 gate( .a(N1863_NOT), .b(EX351), .O(EX352) );
and2 gate( .a(N303), .b(p142), .O(EX353) );
and2 gate( .a(N1863_NOT), .b(EX353), .O(EX354) );
and2 gate( .a(N303_NOT), .b(p143), .O(EX355) );
and2 gate( .a(N1863), .b(EX355), .O(EX356) );
and2 gate( .a(N303), .b(p144), .O(EX357) );
and2 gate( .a(N1863), .b(EX357), .O(EX358) );
or2  gate( .a(EX352), .b(EX354), .O(EX359) );
or2  gate( .a(EX356), .b(EX359), .O(EX360) );
or2  gate( .a(EX358), .b(EX360), .O(N2036) );
and2 gate366( .a(N264), .b(N1864), .O(N2037) );
buf1 gate367( .a(N1667), .O(N2038) );
inv1 gate368( .a(N1667), .O(N2043) );
buf1 gate369( .a(N1670), .O(N2052) );
inv1 gate370( .a(N1670), .O(N2057) );
and3 gate371( .a(N50), .b(N1197), .c(N1869), .O(N2068) );
and3 gate372( .a(N58), .b(N1197), .c(N1874), .O(N2073) );
and3 gate373( .a(N68), .b(N1197), .c(N1879), .O(N2078) );
and3 gate374( .a(N77), .b(N1197), .c(N1884), .O(N2083) );
and3 gate375( .a(N87), .b(N1219), .c(N1889), .O(N2088) );
and3 gate376( .a(N97), .b(N1219), .c(N1894), .O(N2093) );
and3 gate377( .a(N107), .b(N1219), .c(N1899), .O(N2098) );
and3 gate378( .a(N116), .b(N1219), .c(N1904), .O(N2103) );
inv1 gate379( .a(N1562), .O(N2121) );
inv1 gate380( .a(N1562), .O(N2122) );
inv1 gate381( .a(N1562), .O(N2123) );
inv1 gate382( .a(N1562), .O(N2124) );
inv1 gate383( .a(N1562), .O(N2125) );
inv1 gate384( .a(N1562), .O(N2126) );
inv1 gate385( .a(N1562), .O(N2127) );
inv1 gate386( .a(N1562), .O(N2128) );
inv1 gate( .a(N950),.O(N950_NOT) );
inv1 gate( .a(N1939),.O(N1939_NOT));
and2 gate( .a(N950_NOT), .b(p145), .O(EX361) );
and2 gate( .a(N1939_NOT), .b(EX361), .O(EX362) );
and2 gate( .a(N950), .b(p146), .O(EX363) );
and2 gate( .a(N1939_NOT), .b(EX363), .O(EX364) );
and2 gate( .a(N950_NOT), .b(p147), .O(EX365) );
and2 gate( .a(N1939), .b(EX365), .O(EX366) );
and2 gate( .a(N950), .b(p148), .O(EX367) );
and2 gate( .a(N1939), .b(EX367), .O(EX368) );
or2  gate( .a(EX362), .b(EX364), .O(EX369) );
or2  gate( .a(EX366), .b(EX369), .O(EX370) );
or2  gate( .a(EX368), .b(EX370), .O(N2133) );
nand2 gate388( .a(N1478), .b(N1941), .O(N2134) );
nand2 gate389( .a(N1475), .b(N1942), .O(N2135) );
nand2 gate390( .a(N1484), .b(N1943), .O(N2136) );
inv1 gate( .a(N1481),.O(N1481_NOT) );
inv1 gate( .a(N1944),.O(N1944_NOT));
and2 gate( .a(N1481_NOT), .b(p149), .O(EX371) );
and2 gate( .a(N1944_NOT), .b(EX371), .O(EX372) );
and2 gate( .a(N1481), .b(p150), .O(EX373) );
and2 gate( .a(N1944_NOT), .b(EX373), .O(EX374) );
and2 gate( .a(N1481_NOT), .b(p151), .O(EX375) );
and2 gate( .a(N1944), .b(EX375), .O(EX376) );
and2 gate( .a(N1481), .b(p152), .O(EX377) );
and2 gate( .a(N1944), .b(EX377), .O(EX378) );
or2  gate( .a(EX372), .b(EX374), .O(EX379) );
or2  gate( .a(EX376), .b(EX379), .O(EX380) );
or2  gate( .a(EX378), .b(EX380), .O(N2137) );
nand2 gate392( .a(N1490), .b(N1945), .O(N2138) );
inv1 gate( .a(N1487),.O(N1487_NOT) );
inv1 gate( .a(N1946),.O(N1946_NOT));
and2 gate( .a(N1487_NOT), .b(p153), .O(EX381) );
and2 gate( .a(N1946_NOT), .b(EX381), .O(EX382) );
and2 gate( .a(N1487), .b(p154), .O(EX383) );
and2 gate( .a(N1946_NOT), .b(EX383), .O(EX384) );
and2 gate( .a(N1487_NOT), .b(p155), .O(EX385) );
and2 gate( .a(N1946), .b(EX385), .O(EX386) );
and2 gate( .a(N1487), .b(p156), .O(EX387) );
and2 gate( .a(N1946), .b(EX387), .O(EX388) );
or2  gate( .a(EX382), .b(EX384), .O(EX389) );
or2  gate( .a(EX386), .b(EX389), .O(EX390) );
or2  gate( .a(EX388), .b(EX390), .O(N2139) );
inv1 gate394( .a(N1933), .O(N2141) );
inv1 gate395( .a(N1936), .O(N2142) );
inv1 gate396( .a(N1738), .O(N2143) );
and2 gate397( .a(N1738), .b(N1747), .O(N2144) );
inv1 gate398( .a(N1747), .O(N2145) );
nand2 gate399( .a(N1727), .b(N1960), .O(N2146) );
nand2 gate400( .a(N1730), .b(N1961), .O(N2147) );
and4 gate401( .a(N1722), .b(N1267), .c(N665), .d(N58), .O(N2148) );
inv1 gate402( .a(N1738), .O(N2149) );
and2 gate403( .a(N1738), .b(N1747), .O(N2150) );
inv1 gate404( .a(N1747), .O(N2151) );
inv1 gate405( .a(N1738), .O(N2152) );
inv1 gate406( .a(N1747), .O(N2153) );
and2 gate407( .a(N1738), .b(N1747), .O(N2154) );
inv1 gate408( .a(N1738), .O(N2155) );
inv1 gate409( .a(N1747), .O(N2156) );
and2 gate410( .a(N1738), .b(N1747), .O(N2157) );
buf1 gate411( .a(N1761), .O(N2158) );
buf1 gate412( .a(N1761), .O(N2175) );
nand2 gate413( .a(N1764), .b(N1981), .O(N2178) );
nand2 gate414( .a(N1766), .b(N1982), .O(N2179) );
inv1 gate415( .a(N1756), .O(N2180) );
and2 gate416( .a(N1756), .b(N1328), .O(N2181) );
inv1 gate417( .a(N1756), .O(N2183) );
and2 gate418( .a(N1331), .b(N1756), .O(N2184) );
nand2 gate419( .a(N1358), .b(N1812), .O(N2185) );
nand2 gate420( .a(N1358), .b(N1809), .O(N2188) );
inv1 gate( .a(N1353),.O(N1353_NOT) );
inv1 gate( .a(N1812),.O(N1812_NOT));
and2 gate( .a(N1353_NOT), .b(p157), .O(EX391) );
and2 gate( .a(N1812_NOT), .b(EX391), .O(EX392) );
and2 gate( .a(N1353), .b(p158), .O(EX393) );
and2 gate( .a(N1812_NOT), .b(EX393), .O(EX394) );
and2 gate( .a(N1353_NOT), .b(p159), .O(EX395) );
and2 gate( .a(N1812), .b(EX395), .O(EX396) );
and2 gate( .a(N1353), .b(p160), .O(EX397) );
and2 gate( .a(N1812), .b(EX397), .O(EX398) );
or2  gate( .a(EX392), .b(EX394), .O(EX399) );
or2  gate( .a(EX396), .b(EX399), .O(EX400) );
or2  gate( .a(EX398), .b(EX400), .O(N2191) );
nand2 gate422( .a(N1353), .b(N1809), .O(N2194) );
nand2 gate423( .a(N1358), .b(N1806), .O(N2197) );
nand2 gate424( .a(N1358), .b(N1803), .O(N2200) );
nand2 gate425( .a(N1353), .b(N1806), .O(N2203) );
nand2 gate426( .a(N1353), .b(N1803), .O(N2206) );
inv1 gate427( .a(N1815), .O(N2209) );
inv1 gate428( .a(N1818), .O(N2210) );
and2 gate429( .a(N1815), .b(N1818), .O(N2211) );
buf1 gate430( .a(N1821), .O(N2212) );
buf1 gate431( .a(N1821), .O(N2221) );
inv1 gate432( .a(N1833), .O(N2230) );
inv1 gate433( .a(N1833), .O(N2231) );
inv1 gate434( .a(N1833), .O(N2232) );
inv1 gate435( .a(N1833), .O(N2233) );
inv1 gate436( .a(N1824), .O(N2234) );
inv1 gate437( .a(N1824), .O(N2235) );
inv1 gate438( .a(N1824), .O(N2236) );
inv1 gate439( .a(N1824), .O(N2237) );
or3 gate440( .a(N2022), .b(N1643), .c(N2023), .O(N2238) );
or3 gate441( .a(N2024), .b(N1644), .c(N2025), .O(N2239) );
or3 gate442( .a(N2026), .b(N1645), .c(N2027), .O(N2240) );
or3 gate443( .a(N2028), .b(N1646), .c(N2029), .O(N2241) );
or3 gate444( .a(N2030), .b(N1647), .c(N2031), .O(N2242) );
or3 gate445( .a(N2032), .b(N1648), .c(N2033), .O(N2243) );
or3 gate446( .a(N2034), .b(N1649), .c(N2035), .O(N2244) );
or3 gate447( .a(N2036), .b(N1650), .c(N2037), .O(N2245) );
and2 gate448( .a(N1986), .b(N1673), .O(N2270) );
and2 gate449( .a(N1987), .b(N1675), .O(N2277) );
and2 gate450( .a(N1988), .b(N1676), .O(N2282) );
and2 gate451( .a(N1989), .b(N1677), .O(N2287) );
and2 gate452( .a(N1990), .b(N1679), .O(N2294) );
and2 gate453( .a(N1991), .b(N1680), .O(N2299) );
buf1 gate454( .a(N1917), .O(N2304) );
inv1 gate( .a(N1930),.O(N1930_NOT) );
inv1 gate( .a(N350),.O(N350_NOT));
and2 gate( .a(N1930_NOT), .b(p161), .O(EX401) );
and2 gate( .a(N350_NOT), .b(EX401), .O(EX402) );
and2 gate( .a(N1930), .b(p162), .O(EX403) );
and2 gate( .a(N350_NOT), .b(EX403), .O(EX404) );
and2 gate( .a(N1930_NOT), .b(p163), .O(EX405) );
and2 gate( .a(N350), .b(EX405), .O(EX406) );
and2 gate( .a(N1930), .b(p164), .O(EX407) );
and2 gate( .a(N350), .b(EX407), .O(EX408) );
or2  gate( .a(EX402), .b(EX404), .O(EX409) );
or2  gate( .a(EX406), .b(EX409), .O(EX410) );
or2  gate( .a(EX408), .b(EX410), .O(N2307) );
inv1 gate( .a(N1930),.O(N1930_NOT) );
inv1 gate( .a(N350),.O(N350_NOT));
and2 gate( .a(N1930_NOT), .b(p165), .O(EX411) );
and2 gate( .a(N350_NOT), .b(EX411), .O(EX412) );
and2 gate( .a(N1930), .b(p166), .O(EX413) );
and2 gate( .a(N350_NOT), .b(EX413), .O(EX414) );
and2 gate( .a(N1930_NOT), .b(p167), .O(EX415) );
and2 gate( .a(N350), .b(EX415), .O(EX416) );
and2 gate( .a(N1930), .b(p168), .O(EX417) );
and2 gate( .a(N350), .b(EX417), .O(EX418) );
or2  gate( .a(EX412), .b(EX414), .O(EX419) );
or2  gate( .a(EX416), .b(EX419), .O(EX420) );
or2  gate( .a(EX418), .b(EX420), .O(N2310) );
buf1 gate457( .a(N1715), .O(N2313) );
buf1 gate458( .a(N1718), .O(N2316) );
buf1 gate459( .a(N1715), .O(N2319) );
buf1 gate460( .a(N1718), .O(N2322) );
nand2 gate461( .a(N1940), .b(N2133), .O(N2325) );
nand2 gate462( .a(N2134), .b(N2135), .O(N2328) );
nand2 gate463( .a(N2136), .b(N2137), .O(N2331) );
nand2 gate464( .a(N2138), .b(N2139), .O(N2334) );
nand2 gate465( .a(N1936), .b(N2141), .O(N2341) );
inv1 gate( .a(N1933),.O(N1933_NOT) );
inv1 gate( .a(N2142),.O(N2142_NOT));
and2 gate( .a(N1933_NOT), .b(p169), .O(EX421) );
and2 gate( .a(N2142_NOT), .b(EX421), .O(EX422) );
and2 gate( .a(N1933), .b(p170), .O(EX423) );
and2 gate( .a(N2142_NOT), .b(EX423), .O(EX424) );
and2 gate( .a(N1933_NOT), .b(p171), .O(EX425) );
and2 gate( .a(N2142), .b(EX425), .O(EX426) );
and2 gate( .a(N1933), .b(p172), .O(EX427) );
and2 gate( .a(N2142), .b(EX427), .O(EX428) );
or2  gate( .a(EX422), .b(EX424), .O(EX429) );
or2  gate( .a(EX426), .b(EX429), .O(EX430) );
or2  gate( .a(EX428), .b(EX430), .O(N2342) );
and2 gate467( .a(N724), .b(N2144), .O(N2347) );
and3 gate468( .a(N2146), .b(N699), .c(N1726), .O(N2348) );
and2 gate469( .a(N753), .b(N2147), .O(N2349) );
and2 gate470( .a(N2148), .b(N1273), .O(N2350) );
and2 gate471( .a(N736), .b(N2150), .O(N2351) );
and2 gate472( .a(N1735), .b(N2153), .O(N2352) );
inv1 gate( .a(N763),.O(N763_NOT) );
inv1 gate( .a(N2154),.O(N2154_NOT));
and2 gate( .a(N763_NOT), .b(p173), .O(EX431) );
and2 gate( .a(N2154_NOT), .b(EX431), .O(EX432) );
and2 gate( .a(N763), .b(p174), .O(EX433) );
and2 gate( .a(N2154_NOT), .b(EX433), .O(EX434) );
and2 gate( .a(N763_NOT), .b(p175), .O(EX435) );
and2 gate( .a(N2154), .b(EX435), .O(EX436) );
and2 gate( .a(N763), .b(p176), .O(EX437) );
and2 gate( .a(N2154), .b(EX437), .O(EX438) );
or2  gate( .a(EX432), .b(EX434), .O(EX439) );
or2  gate( .a(EX436), .b(EX439), .O(EX440) );
or2  gate( .a(EX438), .b(EX440), .O(N2353) );
inv1 gate( .a(N1725),.O(N1725_NOT) );
inv1 gate( .a(N2156),.O(N2156_NOT));
and2 gate( .a(N1725_NOT), .b(p177), .O(EX441) );
and2 gate( .a(N2156_NOT), .b(EX441), .O(EX442) );
and2 gate( .a(N1725), .b(p178), .O(EX443) );
and2 gate( .a(N2156_NOT), .b(EX443), .O(EX444) );
and2 gate( .a(N1725_NOT), .b(p179), .O(EX445) );
and2 gate( .a(N2156), .b(EX445), .O(EX446) );
and2 gate( .a(N1725), .b(p180), .O(EX447) );
and2 gate( .a(N2156), .b(EX447), .O(EX448) );
or2  gate( .a(EX442), .b(EX444), .O(EX449) );
or2  gate( .a(EX446), .b(EX449), .O(EX450) );
or2  gate( .a(EX448), .b(EX450), .O(N2354) );
and2 gate475( .a(N749), .b(N2157), .O(N2355) );
inv1 gate476( .a(N2178), .O(N2374) );
inv1 gate477( .a(N2179), .O(N2375) );
inv1 gate( .a(N1520),.O(N1520_NOT) );
inv1 gate( .a(N2180),.O(N2180_NOT));
and2 gate( .a(N1520_NOT), .b(p181), .O(EX451) );
and2 gate( .a(N2180_NOT), .b(EX451), .O(EX452) );
and2 gate( .a(N1520), .b(p182), .O(EX453) );
and2 gate( .a(N2180_NOT), .b(EX453), .O(EX454) );
and2 gate( .a(N1520_NOT), .b(p183), .O(EX455) );
and2 gate( .a(N2180), .b(EX455), .O(EX456) );
and2 gate( .a(N1520), .b(p184), .O(EX457) );
and2 gate( .a(N2180), .b(EX457), .O(EX458) );
or2  gate( .a(EX452), .b(EX454), .O(EX459) );
or2  gate( .a(EX456), .b(EX459), .O(EX460) );
or2  gate( .a(EX458), .b(EX460), .O(N2376) );
inv1 gate( .a(N1721),.O(N1721_NOT) );
inv1 gate( .a(N2181),.O(N2181_NOT));
and2 gate( .a(N1721_NOT), .b(p185), .O(EX461) );
and2 gate( .a(N2181_NOT), .b(EX461), .O(EX462) );
and2 gate( .a(N1721), .b(p186), .O(EX463) );
and2 gate( .a(N2181_NOT), .b(EX463), .O(EX464) );
and2 gate( .a(N1721_NOT), .b(p187), .O(EX465) );
and2 gate( .a(N2181), .b(EX465), .O(EX466) );
and2 gate( .a(N1721), .b(p188), .O(EX467) );
and2 gate( .a(N2181), .b(EX467), .O(EX468) );
or2  gate( .a(EX462), .b(EX464), .O(EX469) );
or2  gate( .a(EX466), .b(EX469), .O(EX470) );
or2  gate( .a(EX468), .b(EX470), .O(N2379) );
and2 gate480( .a(N665), .b(N2211), .O(N2398) );
and3 gate481( .a(N2057), .b(N226), .c(N1873), .O(N2417) );
and3 gate482( .a(N2057), .b(N274), .c(N1306), .O(N2418) );
inv1 gate( .a(N2052),.O(N2052_NOT) );
inv1 gate( .a(N2238),.O(N2238_NOT));
and2 gate( .a(N2052_NOT), .b(p189), .O(EX471) );
and2 gate( .a(N2238_NOT), .b(EX471), .O(EX472) );
and2 gate( .a(N2052), .b(p190), .O(EX473) );
and2 gate( .a(N2238_NOT), .b(EX473), .O(EX474) );
and2 gate( .a(N2052_NOT), .b(p191), .O(EX475) );
and2 gate( .a(N2238), .b(EX475), .O(EX476) );
and2 gate( .a(N2052), .b(p192), .O(EX477) );
and2 gate( .a(N2238), .b(EX477), .O(EX478) );
or2  gate( .a(EX472), .b(EX474), .O(EX479) );
or2  gate( .a(EX476), .b(EX479), .O(EX480) );
or2  gate( .a(EX478), .b(EX480), .O(N2419) );
and3 gate484( .a(N2057), .b(N232), .c(N1878), .O(N2420) );
and3 gate485( .a(N2057), .b(N274), .c(N1306), .O(N2421) );
inv1 gate( .a(N2052),.O(N2052_NOT) );
inv1 gate( .a(N2239),.O(N2239_NOT));
and2 gate( .a(N2052_NOT), .b(p193), .O(EX481) );
and2 gate( .a(N2239_NOT), .b(EX481), .O(EX482) );
and2 gate( .a(N2052), .b(p194), .O(EX483) );
and2 gate( .a(N2239_NOT), .b(EX483), .O(EX484) );
and2 gate( .a(N2052_NOT), .b(p195), .O(EX485) );
and2 gate( .a(N2239), .b(EX485), .O(EX486) );
and2 gate( .a(N2052), .b(p196), .O(EX487) );
and2 gate( .a(N2239), .b(EX487), .O(EX488) );
or2  gate( .a(EX482), .b(EX484), .O(EX489) );
or2  gate( .a(EX486), .b(EX489), .O(EX490) );
or2  gate( .a(EX488), .b(EX490), .O(N2422) );
and3 gate487( .a(N2057), .b(N238), .c(N1883), .O(N2425) );
and3 gate488( .a(N2057), .b(N274), .c(N1306), .O(N2426) );
and2 gate489( .a(N2052), .b(N2240), .O(N2427) );
and3 gate490( .a(N2057), .b(N244), .c(N1888), .O(N2430) );
and3 gate491( .a(N2057), .b(N274), .c(N1306), .O(N2431) );
and2 gate492( .a(N2052), .b(N2241), .O(N2432) );
and3 gate493( .a(N2043), .b(N250), .c(N1893), .O(N2435) );
and3 gate494( .a(N2043), .b(N274), .c(N1322), .O(N2436) );
inv1 gate( .a(N2038),.O(N2038_NOT) );
inv1 gate( .a(N2242),.O(N2242_NOT));
and2 gate( .a(N2038_NOT), .b(p197), .O(EX491) );
and2 gate( .a(N2242_NOT), .b(EX491), .O(EX492) );
and2 gate( .a(N2038), .b(p198), .O(EX493) );
and2 gate( .a(N2242_NOT), .b(EX493), .O(EX494) );
and2 gate( .a(N2038_NOT), .b(p199), .O(EX495) );
and2 gate( .a(N2242), .b(EX495), .O(EX496) );
and2 gate( .a(N2038), .b(p200), .O(EX497) );
and2 gate( .a(N2242), .b(EX497), .O(EX498) );
or2  gate( .a(EX492), .b(EX494), .O(EX499) );
or2  gate( .a(EX496), .b(EX499), .O(EX500) );
or2  gate( .a(EX498), .b(EX500), .O(N2437) );
and3 gate496( .a(N2043), .b(N257), .c(N1898), .O(N2438) );
and3 gate497( .a(N2043), .b(N274), .c(N1315), .O(N2439) );
and2 gate498( .a(N2038), .b(N2243), .O(N2440) );
and3 gate499( .a(N2043), .b(N264), .c(N1903), .O(N2443) );
and3 gate500( .a(N2043), .b(N274), .c(N1315), .O(N2444) );
and2 gate501( .a(N2038), .b(N2244), .O(N2445) );
and3 gate502( .a(N2043), .b(N270), .c(N1908), .O(N2448) );
and3 gate503( .a(N2043), .b(N274), .c(N1315), .O(N2449) );
and2 gate504( .a(N2038), .b(N2245), .O(N2450) );
inv1 gate505( .a(N2313), .O(N2467) );
inv1 gate506( .a(N2316), .O(N2468) );
inv1 gate507( .a(N2319), .O(N2469) );
inv1 gate508( .a(N2322), .O(N2470) );
nand2 gate509( .a(N2341), .b(N2342), .O(N2471) );
inv1 gate510( .a(N2325), .O(N2474) );
inv1 gate511( .a(N2328), .O(N2475) );
inv1 gate512( .a(N2331), .O(N2476) );
inv1 gate513( .a(N2334), .O(N2477) );
inv1 gate( .a(N2348),.O(N2348_NOT) );
inv1 gate( .a(N1729),.O(N1729_NOT));
and2 gate( .a(N2348_NOT), .b(p201), .O(EX501) );
and2 gate( .a(N1729_NOT), .b(EX501), .O(EX502) );
and2 gate( .a(N2348), .b(p202), .O(EX503) );
and2 gate( .a(N1729_NOT), .b(EX503), .O(EX504) );
and2 gate( .a(N2348_NOT), .b(p203), .O(EX505) );
and2 gate( .a(N1729), .b(EX505), .O(EX506) );
and2 gate( .a(N2348), .b(p204), .O(EX507) );
and2 gate( .a(N1729), .b(EX507), .O(EX508) );
or2  gate( .a(EX502), .b(EX504), .O(EX509) );
or2  gate( .a(EX506), .b(EX509), .O(EX510) );
or2  gate( .a(EX508), .b(EX510), .O(N2478) );
inv1 gate515( .a(N2175), .O(N2481) );
inv1 gate( .a(N2175),.O(N2175_NOT) );
inv1 gate( .a(N1334),.O(N1334_NOT));
and2 gate( .a(N2175_NOT), .b(p205), .O(EX511) );
and2 gate( .a(N1334_NOT), .b(EX511), .O(EX512) );
and2 gate( .a(N2175), .b(p206), .O(EX513) );
and2 gate( .a(N1334_NOT), .b(EX513), .O(EX514) );
and2 gate( .a(N2175_NOT), .b(p207), .O(EX515) );
and2 gate( .a(N1334), .b(EX515), .O(EX516) );
and2 gate( .a(N2175), .b(p208), .O(EX517) );
and2 gate( .a(N1334), .b(EX517), .O(EX518) );
or2  gate( .a(EX512), .b(EX514), .O(EX519) );
or2  gate( .a(EX516), .b(EX519), .O(EX520) );
or2  gate( .a(EX518), .b(EX520), .O(N2482) );
inv1 gate( .a(N2349),.O(N2349_NOT) );
inv1 gate( .a(N2183),.O(N2183_NOT));
and2 gate( .a(N2349_NOT), .b(p209), .O(EX521) );
and2 gate( .a(N2183_NOT), .b(EX521), .O(EX522) );
and2 gate( .a(N2349), .b(p210), .O(EX523) );
and2 gate( .a(N2183_NOT), .b(EX523), .O(EX524) );
and2 gate( .a(N2349_NOT), .b(p211), .O(EX525) );
and2 gate( .a(N2183), .b(EX525), .O(EX526) );
and2 gate( .a(N2349), .b(p212), .O(EX527) );
and2 gate( .a(N2183), .b(EX527), .O(EX528) );
or2  gate( .a(EX522), .b(EX524), .O(EX529) );
or2  gate( .a(EX526), .b(EX529), .O(EX530) );
or2  gate( .a(EX528), .b(EX530), .O(N2483) );
and2 gate518( .a(N2374), .b(N1346), .O(N2486) );
and2 gate519( .a(N2375), .b(N1350), .O(N2487) );
buf1 gate520( .a(N2185), .O(N2488) );
buf1 gate521( .a(N2188), .O(N2497) );
buf1 gate522( .a(N2191), .O(N2506) );
buf1 gate523( .a(N2194), .O(N2515) );
buf1 gate524( .a(N2197), .O(N2524) );
buf1 gate525( .a(N2200), .O(N2533) );
buf1 gate526( .a(N2203), .O(N2542) );
buf1 gate527( .a(N2206), .O(N2551) );
buf1 gate528( .a(N2185), .O(N2560) );
buf1 gate529( .a(N2188), .O(N2569) );
buf1 gate530( .a(N2191), .O(N2578) );
buf1 gate531( .a(N2194), .O(N2587) );
buf1 gate532( .a(N2197), .O(N2596) );
buf1 gate533( .a(N2200), .O(N2605) );
buf1 gate534( .a(N2203), .O(N2614) );
buf1 gate535( .a(N2206), .O(N2623) );
inv1 gate536( .a(N2212), .O(N2632) );
and2 gate537( .a(N2212), .b(N1833), .O(N2633) );
inv1 gate538( .a(N2212), .O(N2634) );
and2 gate539( .a(N2212), .b(N1833), .O(N2635) );
inv1 gate540( .a(N2212), .O(N2636) );
inv1 gate( .a(N2212),.O(N2212_NOT) );
inv1 gate( .a(N1833),.O(N1833_NOT));
and2 gate( .a(N2212_NOT), .b(p213), .O(EX531) );
and2 gate( .a(N1833_NOT), .b(EX531), .O(EX532) );
and2 gate( .a(N2212), .b(p214), .O(EX533) );
and2 gate( .a(N1833_NOT), .b(EX533), .O(EX534) );
and2 gate( .a(N2212_NOT), .b(p215), .O(EX535) );
and2 gate( .a(N1833), .b(EX535), .O(EX536) );
and2 gate( .a(N2212), .b(p216), .O(EX537) );
and2 gate( .a(N1833), .b(EX537), .O(EX538) );
or2  gate( .a(EX532), .b(EX534), .O(EX539) );
or2  gate( .a(EX536), .b(EX539), .O(EX540) );
or2  gate( .a(EX538), .b(EX540), .O(N2637) );
inv1 gate542( .a(N2212), .O(N2638) );
and2 gate543( .a(N2212), .b(N1833), .O(N2639) );
inv1 gate544( .a(N2221), .O(N2640) );
and2 gate545( .a(N2221), .b(N1824), .O(N2641) );
inv1 gate546( .a(N2221), .O(N2642) );
and2 gate547( .a(N2221), .b(N1824), .O(N2643) );
inv1 gate548( .a(N2221), .O(N2644) );
and2 gate549( .a(N2221), .b(N1824), .O(N2645) );
inv1 gate550( .a(N2221), .O(N2646) );
and2 gate551( .a(N2221), .b(N1824), .O(N2647) );
or3 gate552( .a(N2270), .b(N1870), .c(N2068), .O(N2648) );
nor3 gate553( .a(N2270), .b(N1870), .c(N2068), .O(N2652) );
or3 gate554( .a(N2417), .b(N2418), .c(N2419), .O(N2656) );
or3 gate555( .a(N2420), .b(N2421), .c(N2422), .O(N2659) );
or3 gate556( .a(N2277), .b(N1880), .c(N2078), .O(N2662) );
nor3 gate557( .a(N2277), .b(N1880), .c(N2078), .O(N2666) );
or3 gate558( .a(N2425), .b(N2426), .c(N2427), .O(N2670) );
or3 gate559( .a(N2282), .b(N1885), .c(N2083), .O(N2673) );
nor3 gate560( .a(N2282), .b(N1885), .c(N2083), .O(N2677) );
or3 gate561( .a(N2430), .b(N2431), .c(N2432), .O(N2681) );
or3 gate562( .a(N2287), .b(N1890), .c(N2088), .O(N2684) );
nor3 gate563( .a(N2287), .b(N1890), .c(N2088), .O(N2688) );
or3 gate564( .a(N2435), .b(N2436), .c(N2437), .O(N2692) );
or3 gate565( .a(N2438), .b(N2439), .c(N2440), .O(N2697) );
or3 gate566( .a(N2294), .b(N1900), .c(N2098), .O(N2702) );
nor3 gate567( .a(N2294), .b(N1900), .c(N2098), .O(N2706) );
or3 gate568( .a(N2443), .b(N2444), .c(N2445), .O(N2710) );
or3 gate569( .a(N2299), .b(N1905), .c(N2103), .O(N2715) );
nor3 gate570( .a(N2299), .b(N1905), .c(N2103), .O(N2719) );
or3 gate571( .a(N2448), .b(N2449), .c(N2450), .O(N2723) );
inv1 gate572( .a(N2304), .O(N2728) );
inv1 gate573( .a(N2158), .O(N2729) );
inv1 gate( .a(N1562),.O(N1562_NOT) );
inv1 gate( .a(N2158),.O(N2158_NOT));
and2 gate( .a(N1562_NOT), .b(p217), .O(EX541) );
and2 gate( .a(N2158_NOT), .b(EX541), .O(EX542) );
and2 gate( .a(N1562), .b(p218), .O(EX543) );
and2 gate( .a(N2158_NOT), .b(EX543), .O(EX544) );
and2 gate( .a(N1562_NOT), .b(p219), .O(EX545) );
and2 gate( .a(N2158), .b(EX545), .O(EX546) );
and2 gate( .a(N1562), .b(p220), .O(EX547) );
and2 gate( .a(N2158), .b(EX547), .O(EX548) );
or2  gate( .a(EX542), .b(EX544), .O(EX549) );
or2  gate( .a(EX546), .b(EX549), .O(EX550) );
or2  gate( .a(EX548), .b(EX550), .O(N2730) );
inv1 gate575( .a(N2158), .O(N2731) );
and2 gate576( .a(N1562), .b(N2158), .O(N2732) );
inv1 gate577( .a(N2158), .O(N2733) );
and2 gate578( .a(N1562), .b(N2158), .O(N2734) );
inv1 gate579( .a(N2158), .O(N2735) );
and2 gate580( .a(N1562), .b(N2158), .O(N2736) );
inv1 gate581( .a(N2158), .O(N2737) );
and2 gate582( .a(N1562), .b(N2158), .O(N2738) );
inv1 gate583( .a(N2158), .O(N2739) );
and2 gate584( .a(N1562), .b(N2158), .O(N2740) );
inv1 gate585( .a(N2158), .O(N2741) );
inv1 gate( .a(N1562),.O(N1562_NOT) );
inv1 gate( .a(N2158),.O(N2158_NOT));
and2 gate( .a(N1562_NOT), .b(p221), .O(EX551) );
and2 gate( .a(N2158_NOT), .b(EX551), .O(EX552) );
and2 gate( .a(N1562), .b(p222), .O(EX553) );
and2 gate( .a(N2158_NOT), .b(EX553), .O(EX554) );
and2 gate( .a(N1562_NOT), .b(p223), .O(EX555) );
and2 gate( .a(N2158), .b(EX555), .O(EX556) );
and2 gate( .a(N1562), .b(p224), .O(EX557) );
and2 gate( .a(N2158), .b(EX557), .O(EX558) );
or2  gate( .a(EX552), .b(EX554), .O(EX559) );
or2  gate( .a(EX556), .b(EX559), .O(EX560) );
or2  gate( .a(EX558), .b(EX560), .O(N2742) );
inv1 gate587( .a(N2158), .O(N2743) );
and2 gate588( .a(N1562), .b(N2158), .O(N2744) );
or3 gate589( .a(N2376), .b(N1983), .c(N2379), .O(N2745) );
nor3 gate590( .a(N2376), .b(N1983), .c(N2379), .O(N2746) );
inv1 gate( .a(N2316),.O(N2316_NOT) );
inv1 gate( .a(N2467),.O(N2467_NOT));
and2 gate( .a(N2316_NOT), .b(p225), .O(EX561) );
and2 gate( .a(N2467_NOT), .b(EX561), .O(EX562) );
and2 gate( .a(N2316), .b(p226), .O(EX563) );
and2 gate( .a(N2467_NOT), .b(EX563), .O(EX564) );
and2 gate( .a(N2316_NOT), .b(p227), .O(EX565) );
and2 gate( .a(N2467), .b(EX565), .O(EX566) );
and2 gate( .a(N2316), .b(p228), .O(EX567) );
and2 gate( .a(N2467), .b(EX567), .O(EX568) );
or2  gate( .a(EX562), .b(EX564), .O(EX569) );
or2  gate( .a(EX566), .b(EX569), .O(EX570) );
or2  gate( .a(EX568), .b(EX570), .O(N2748) );
nand2 gate592( .a(N2313), .b(N2468), .O(N2749) );
nand2 gate593( .a(N2322), .b(N2469), .O(N2750) );
nand2 gate594( .a(N2319), .b(N2470), .O(N2751) );
nand2 gate595( .a(N2328), .b(N2474), .O(N2754) );
inv1 gate( .a(N2325),.O(N2325_NOT) );
inv1 gate( .a(N2475),.O(N2475_NOT));
and2 gate( .a(N2325_NOT), .b(p229), .O(EX571) );
and2 gate( .a(N2475_NOT), .b(EX571), .O(EX572) );
and2 gate( .a(N2325), .b(p230), .O(EX573) );
and2 gate( .a(N2475_NOT), .b(EX573), .O(EX574) );
and2 gate( .a(N2325_NOT), .b(p231), .O(EX575) );
and2 gate( .a(N2475), .b(EX575), .O(EX576) );
and2 gate( .a(N2325), .b(p232), .O(EX577) );
and2 gate( .a(N2475), .b(EX577), .O(EX578) );
or2  gate( .a(EX572), .b(EX574), .O(EX579) );
or2  gate( .a(EX576), .b(EX579), .O(EX580) );
or2  gate( .a(EX578), .b(EX580), .O(N2755) );
nand2 gate597( .a(N2334), .b(N2476), .O(N2756) );
nand2 gate598( .a(N2331), .b(N2477), .O(N2757) );
inv1 gate( .a(N1520),.O(N1520_NOT) );
inv1 gate( .a(N2481),.O(N2481_NOT));
and2 gate( .a(N1520_NOT), .b(p233), .O(EX581) );
and2 gate( .a(N2481_NOT), .b(EX581), .O(EX582) );
and2 gate( .a(N1520), .b(p234), .O(EX583) );
and2 gate( .a(N2481_NOT), .b(EX583), .O(EX584) );
and2 gate( .a(N1520_NOT), .b(p235), .O(EX585) );
and2 gate( .a(N2481), .b(EX585), .O(EX586) );
and2 gate( .a(N1520), .b(p236), .O(EX587) );
and2 gate( .a(N2481), .b(EX587), .O(EX588) );
or2  gate( .a(EX582), .b(EX584), .O(EX589) );
or2  gate( .a(EX586), .b(EX589), .O(EX590) );
or2  gate( .a(EX588), .b(EX590), .O(N2758) );
inv1 gate( .a(N1722),.O(N1722_NOT) );
inv1 gate( .a(N2482),.O(N2482_NOT));
and2 gate( .a(N1722_NOT), .b(p237), .O(EX591) );
and2 gate( .a(N2482_NOT), .b(EX591), .O(EX592) );
and2 gate( .a(N1722), .b(p238), .O(EX593) );
and2 gate( .a(N2482_NOT), .b(EX593), .O(EX594) );
and2 gate( .a(N1722_NOT), .b(p239), .O(EX595) );
and2 gate( .a(N2482), .b(EX595), .O(EX596) );
and2 gate( .a(N1722), .b(p240), .O(EX597) );
and2 gate( .a(N2482), .b(EX597), .O(EX598) );
or2  gate( .a(EX592), .b(EX594), .O(EX599) );
or2  gate( .a(EX596), .b(EX599), .O(EX600) );
or2  gate( .a(EX598), .b(EX600), .O(N2761) );
and2 gate601( .a(N2478), .b(N1770), .O(N2764) );
or3 gate602( .a(N2486), .b(N1789), .c(N1790), .O(N2768) );
or3 gate603( .a(N2487), .b(N1797), .c(N1798), .O(N2769) );
inv1 gate( .a(N665),.O(N665_NOT) );
inv1 gate( .a(N2633),.O(N2633_NOT));
and2 gate( .a(N665_NOT), .b(p241), .O(EX601) );
and2 gate( .a(N2633_NOT), .b(EX601), .O(EX602) );
and2 gate( .a(N665), .b(p242), .O(EX603) );
and2 gate( .a(N2633_NOT), .b(EX603), .O(EX604) );
and2 gate( .a(N665_NOT), .b(p243), .O(EX605) );
and2 gate( .a(N2633), .b(EX605), .O(EX606) );
and2 gate( .a(N665), .b(p244), .O(EX607) );
and2 gate( .a(N2633), .b(EX607), .O(EX608) );
or2  gate( .a(EX602), .b(EX604), .O(EX609) );
or2  gate( .a(EX606), .b(EX609), .O(EX610) );
or2  gate( .a(EX608), .b(EX610), .O(N2898) );
and2 gate605( .a(N679), .b(N2635), .O(N2899) );
and2 gate606( .a(N686), .b(N2637), .O(N2900) );
and2 gate607( .a(N702), .b(N2639), .O(N2901) );
inv1 gate608( .a(N2746), .O(N2962) );
nand2 gate609( .a(N2748), .b(N2749), .O(N2966) );
nand2 gate610( .a(N2750), .b(N2751), .O(N2967) );
buf1 gate611( .a(N2471), .O(N2970) );
nand2 gate612( .a(N2754), .b(N2755), .O(N2973) );
nand2 gate613( .a(N2756), .b(N2757), .O(N2977) );
and2 gate614( .a(N2471), .b(N2143), .O(N2980) );
inv1 gate615( .a(N2488), .O(N2984) );
inv1 gate616( .a(N2497), .O(N2985) );
inv1 gate617( .a(N2506), .O(N2986) );
inv1 gate618( .a(N2515), .O(N2987) );
inv1 gate619( .a(N2524), .O(N2988) );
inv1 gate620( .a(N2533), .O(N2989) );
inv1 gate621( .a(N2542), .O(N2990) );
inv1 gate622( .a(N2551), .O(N2991) );
inv1 gate623( .a(N2488), .O(N2992) );
inv1 gate624( .a(N2497), .O(N2993) );
inv1 gate625( .a(N2506), .O(N2994) );
inv1 gate626( .a(N2515), .O(N2995) );
inv1 gate627( .a(N2524), .O(N2996) );
inv1 gate628( .a(N2533), .O(N2997) );
inv1 gate629( .a(N2542), .O(N2998) );
inv1 gate630( .a(N2551), .O(N2999) );
inv1 gate631( .a(N2488), .O(N3000) );
inv1 gate632( .a(N2497), .O(N3001) );
inv1 gate633( .a(N2506), .O(N3002) );
inv1 gate634( .a(N2515), .O(N3003) );
inv1 gate635( .a(N2524), .O(N3004) );
inv1 gate636( .a(N2533), .O(N3005) );
inv1 gate637( .a(N2542), .O(N3006) );
inv1 gate638( .a(N2551), .O(N3007) );
inv1 gate639( .a(N2488), .O(N3008) );
inv1 gate640( .a(N2497), .O(N3009) );
inv1 gate641( .a(N2506), .O(N3010) );
inv1 gate642( .a(N2515), .O(N3011) );
inv1 gate643( .a(N2524), .O(N3012) );
inv1 gate644( .a(N2533), .O(N3013) );
inv1 gate645( .a(N2542), .O(N3014) );
inv1 gate646( .a(N2551), .O(N3015) );
inv1 gate647( .a(N2488), .O(N3016) );
inv1 gate648( .a(N2497), .O(N3017) );
inv1 gate649( .a(N2506), .O(N3018) );
inv1 gate650( .a(N2515), .O(N3019) );
inv1 gate651( .a(N2524), .O(N3020) );
inv1 gate652( .a(N2533), .O(N3021) );
inv1 gate653( .a(N2542), .O(N3022) );
inv1 gate654( .a(N2551), .O(N3023) );
inv1 gate655( .a(N2488), .O(N3024) );
inv1 gate656( .a(N2497), .O(N3025) );
inv1 gate657( .a(N2506), .O(N3026) );
inv1 gate658( .a(N2515), .O(N3027) );
inv1 gate659( .a(N2524), .O(N3028) );
inv1 gate660( .a(N2533), .O(N3029) );
inv1 gate661( .a(N2542), .O(N3030) );
inv1 gate662( .a(N2551), .O(N3031) );
inv1 gate663( .a(N2488), .O(N3032) );
inv1 gate664( .a(N2497), .O(N3033) );
inv1 gate665( .a(N2506), .O(N3034) );
inv1 gate666( .a(N2515), .O(N3035) );
inv1 gate667( .a(N2524), .O(N3036) );
inv1 gate668( .a(N2533), .O(N3037) );
inv1 gate669( .a(N2542), .O(N3038) );
inv1 gate670( .a(N2551), .O(N3039) );
inv1 gate671( .a(N2488), .O(N3040) );
inv1 gate672( .a(N2497), .O(N3041) );
inv1 gate673( .a(N2506), .O(N3042) );
inv1 gate674( .a(N2515), .O(N3043) );
inv1 gate675( .a(N2524), .O(N3044) );
inv1 gate676( .a(N2533), .O(N3045) );
inv1 gate677( .a(N2542), .O(N3046) );
inv1 gate678( .a(N2551), .O(N3047) );
inv1 gate679( .a(N2560), .O(N3048) );
inv1 gate680( .a(N2569), .O(N3049) );
inv1 gate681( .a(N2578), .O(N3050) );
inv1 gate682( .a(N2587), .O(N3051) );
inv1 gate683( .a(N2596), .O(N3052) );
inv1 gate684( .a(N2605), .O(N3053) );
inv1 gate685( .a(N2614), .O(N3054) );
inv1 gate686( .a(N2623), .O(N3055) );
inv1 gate687( .a(N2560), .O(N3056) );
inv1 gate688( .a(N2569), .O(N3057) );
inv1 gate689( .a(N2578), .O(N3058) );
inv1 gate690( .a(N2587), .O(N3059) );
inv1 gate691( .a(N2596), .O(N3060) );
inv1 gate692( .a(N2605), .O(N3061) );
inv1 gate693( .a(N2614), .O(N3062) );
inv1 gate694( .a(N2623), .O(N3063) );
inv1 gate695( .a(N2560), .O(N3064) );
inv1 gate696( .a(N2569), .O(N3065) );
inv1 gate697( .a(N2578), .O(N3066) );
inv1 gate698( .a(N2587), .O(N3067) );
inv1 gate699( .a(N2596), .O(N3068) );
inv1 gate700( .a(N2605), .O(N3069) );
inv1 gate701( .a(N2614), .O(N3070) );
inv1 gate702( .a(N2623), .O(N3071) );
inv1 gate703( .a(N2560), .O(N3072) );
inv1 gate704( .a(N2569), .O(N3073) );
inv1 gate705( .a(N2578), .O(N3074) );
inv1 gate706( .a(N2587), .O(N3075) );
inv1 gate707( .a(N2596), .O(N3076) );
inv1 gate708( .a(N2605), .O(N3077) );
inv1 gate709( .a(N2614), .O(N3078) );
inv1 gate710( .a(N2623), .O(N3079) );
inv1 gate711( .a(N2560), .O(N3080) );
inv1 gate712( .a(N2569), .O(N3081) );
inv1 gate713( .a(N2578), .O(N3082) );
inv1 gate714( .a(N2587), .O(N3083) );
inv1 gate715( .a(N2596), .O(N3084) );
inv1 gate716( .a(N2605), .O(N3085) );
inv1 gate717( .a(N2614), .O(N3086) );
inv1 gate718( .a(N2623), .O(N3087) );
inv1 gate719( .a(N2560), .O(N3088) );
inv1 gate720( .a(N2569), .O(N3089) );
inv1 gate721( .a(N2578), .O(N3090) );
inv1 gate722( .a(N2587), .O(N3091) );
inv1 gate723( .a(N2596), .O(N3092) );
inv1 gate724( .a(N2605), .O(N3093) );
inv1 gate725( .a(N2614), .O(N3094) );
inv1 gate726( .a(N2623), .O(N3095) );
inv1 gate727( .a(N2560), .O(N3096) );
inv1 gate728( .a(N2569), .O(N3097) );
inv1 gate729( .a(N2578), .O(N3098) );
inv1 gate730( .a(N2587), .O(N3099) );
inv1 gate731( .a(N2596), .O(N3100) );
inv1 gate732( .a(N2605), .O(N3101) );
inv1 gate733( .a(N2614), .O(N3102) );
inv1 gate734( .a(N2623), .O(N3103) );
inv1 gate735( .a(N2560), .O(N3104) );
inv1 gate736( .a(N2569), .O(N3105) );
inv1 gate737( .a(N2578), .O(N3106) );
inv1 gate738( .a(N2587), .O(N3107) );
inv1 gate739( .a(N2596), .O(N3108) );
inv1 gate740( .a(N2605), .O(N3109) );
inv1 gate741( .a(N2614), .O(N3110) );
inv1 gate742( .a(N2623), .O(N3111) );
buf1 gate743( .a(N2656), .O(N3112) );
inv1 gate744( .a(N2656), .O(N3115) );
inv1 gate745( .a(N2652), .O(N3118) );
inv1 gate( .a(N2768),.O(N2768_NOT) );
inv1 gate( .a(N1674),.O(N1674_NOT));
and2 gate( .a(N2768_NOT), .b(p245), .O(EX611) );
and2 gate( .a(N1674_NOT), .b(EX611), .O(EX612) );
and2 gate( .a(N2768), .b(p246), .O(EX613) );
and2 gate( .a(N1674_NOT), .b(EX613), .O(EX614) );
and2 gate( .a(N2768_NOT), .b(p247), .O(EX615) );
and2 gate( .a(N1674), .b(EX615), .O(EX616) );
and2 gate( .a(N2768), .b(p248), .O(EX617) );
and2 gate( .a(N1674), .b(EX617), .O(EX618) );
or2  gate( .a(EX612), .b(EX614), .O(EX619) );
or2  gate( .a(EX616), .b(EX619), .O(EX620) );
or2  gate( .a(EX618), .b(EX620), .O(N3119) );
buf1 gate747( .a(N2659), .O(N3122) );
inv1 gate748( .a(N2659), .O(N3125) );
buf1 gate749( .a(N2670), .O(N3128) );
inv1 gate750( .a(N2670), .O(N3131) );
inv1 gate751( .a(N2666), .O(N3134) );
buf1 gate752( .a(N2681), .O(N3135) );
inv1 gate753( .a(N2681), .O(N3138) );
inv1 gate754( .a(N2677), .O(N3141) );
buf1 gate755( .a(N2692), .O(N3142) );
inv1 gate756( .a(N2692), .O(N3145) );
inv1 gate757( .a(N2688), .O(N3148) );
and2 gate758( .a(N2769), .b(N1678), .O(N3149) );
buf1 gate759( .a(N2697), .O(N3152) );
inv1 gate760( .a(N2697), .O(N3155) );
buf1 gate761( .a(N2710), .O(N3158) );
inv1 gate762( .a(N2710), .O(N3161) );
inv1 gate763( .a(N2706), .O(N3164) );
buf1 gate764( .a(N2723), .O(N3165) );
inv1 gate765( .a(N2723), .O(N3168) );
inv1 gate766( .a(N2719), .O(N3171) );
and2 gate767( .a(N1909), .b(N2648), .O(N3172) );
and2 gate768( .a(N1913), .b(N2662), .O(N3175) );
inv1 gate( .a(N1913),.O(N1913_NOT) );
inv1 gate( .a(N2673),.O(N2673_NOT));
and2 gate( .a(N1913_NOT), .b(p249), .O(EX621) );
and2 gate( .a(N2673_NOT), .b(EX621), .O(EX622) );
and2 gate( .a(N1913), .b(p250), .O(EX623) );
and2 gate( .a(N2673_NOT), .b(EX623), .O(EX624) );
and2 gate( .a(N1913_NOT), .b(p251), .O(EX625) );
and2 gate( .a(N2673), .b(EX625), .O(EX626) );
and2 gate( .a(N1913), .b(p252), .O(EX627) );
and2 gate( .a(N2673), .b(EX627), .O(EX628) );
or2  gate( .a(EX622), .b(EX624), .O(EX629) );
or2  gate( .a(EX626), .b(EX629), .O(EX630) );
or2  gate( .a(EX628), .b(EX630), .O(N3178) );
and2 gate770( .a(N1913), .b(N2684), .O(N3181) );
and2 gate771( .a(N1922), .b(N2702), .O(N3184) );
inv1 gate( .a(N1922),.O(N1922_NOT) );
inv1 gate( .a(N2715),.O(N2715_NOT));
and2 gate( .a(N1922_NOT), .b(p253), .O(EX631) );
and2 gate( .a(N2715_NOT), .b(EX631), .O(EX632) );
and2 gate( .a(N1922), .b(p254), .O(EX633) );
and2 gate( .a(N2715_NOT), .b(EX633), .O(EX634) );
and2 gate( .a(N1922_NOT), .b(p255), .O(EX635) );
and2 gate( .a(N2715), .b(EX635), .O(EX636) );
and2 gate( .a(N1922), .b(p256), .O(EX637) );
and2 gate( .a(N2715), .b(EX637), .O(EX638) );
or2  gate( .a(EX632), .b(EX634), .O(EX639) );
or2  gate( .a(EX636), .b(EX639), .O(EX640) );
or2  gate( .a(EX638), .b(EX640), .O(N3187) );
inv1 gate773( .a(N2692), .O(N3190) );
inv1 gate774( .a(N2697), .O(N3191) );
inv1 gate775( .a(N2710), .O(N3192) );
inv1 gate776( .a(N2723), .O(N3193) );
and5 gate777( .a(N2692), .b(N2697), .c(N2710), .d(N2723), .e(N1459), .O(N3194) );
nand2 gate778( .a(N2745), .b(N2962), .O(N3195) );
inv1 gate779( .a(N2966), .O(N3196) );
or3 gate780( .a(N2980), .b(N2145), .c(N2347), .O(N3206) );
and2 gate781( .a(N124), .b(N2984), .O(N3207) );
inv1 gate( .a(N159),.O(N159_NOT) );
inv1 gate( .a(N2985),.O(N2985_NOT));
and2 gate( .a(N159_NOT), .b(p257), .O(EX641) );
and2 gate( .a(N2985_NOT), .b(EX641), .O(EX642) );
and2 gate( .a(N159), .b(p258), .O(EX643) );
and2 gate( .a(N2985_NOT), .b(EX643), .O(EX644) );
and2 gate( .a(N159_NOT), .b(p259), .O(EX645) );
and2 gate( .a(N2985), .b(EX645), .O(EX646) );
and2 gate( .a(N159), .b(p260), .O(EX647) );
and2 gate( .a(N2985), .b(EX647), .O(EX648) );
or2  gate( .a(EX642), .b(EX644), .O(EX649) );
or2  gate( .a(EX646), .b(EX649), .O(EX650) );
or2  gate( .a(EX648), .b(EX650), .O(N3208) );
inv1 gate( .a(N150),.O(N150_NOT) );
inv1 gate( .a(N2986),.O(N2986_NOT));
and2 gate( .a(N150_NOT), .b(p261), .O(EX651) );
and2 gate( .a(N2986_NOT), .b(EX651), .O(EX652) );
and2 gate( .a(N150), .b(p262), .O(EX653) );
and2 gate( .a(N2986_NOT), .b(EX653), .O(EX654) );
and2 gate( .a(N150_NOT), .b(p263), .O(EX655) );
and2 gate( .a(N2986), .b(EX655), .O(EX656) );
and2 gate( .a(N150), .b(p264), .O(EX657) );
and2 gate( .a(N2986), .b(EX657), .O(EX658) );
or2  gate( .a(EX652), .b(EX654), .O(EX659) );
or2  gate( .a(EX656), .b(EX659), .O(EX660) );
or2  gate( .a(EX658), .b(EX660), .O(N3209) );
inv1 gate( .a(N143),.O(N143_NOT) );
inv1 gate( .a(N2987),.O(N2987_NOT));
and2 gate( .a(N143_NOT), .b(p265), .O(EX661) );
and2 gate( .a(N2987_NOT), .b(EX661), .O(EX662) );
and2 gate( .a(N143), .b(p266), .O(EX663) );
and2 gate( .a(N2987_NOT), .b(EX663), .O(EX664) );
and2 gate( .a(N143_NOT), .b(p267), .O(EX665) );
and2 gate( .a(N2987), .b(EX665), .O(EX666) );
and2 gate( .a(N143), .b(p268), .O(EX667) );
and2 gate( .a(N2987), .b(EX667), .O(EX668) );
or2  gate( .a(EX662), .b(EX664), .O(EX669) );
or2  gate( .a(EX666), .b(EX669), .O(EX670) );
or2  gate( .a(EX668), .b(EX670), .O(N3210) );
and2 gate785( .a(N137), .b(N2988), .O(N3211) );
inv1 gate( .a(N132),.O(N132_NOT) );
inv1 gate( .a(N2989),.O(N2989_NOT));
and2 gate( .a(N132_NOT), .b(p269), .O(EX671) );
and2 gate( .a(N2989_NOT), .b(EX671), .O(EX672) );
and2 gate( .a(N132), .b(p270), .O(EX673) );
and2 gate( .a(N2989_NOT), .b(EX673), .O(EX674) );
and2 gate( .a(N132_NOT), .b(p271), .O(EX675) );
and2 gate( .a(N2989), .b(EX675), .O(EX676) );
and2 gate( .a(N132), .b(p272), .O(EX677) );
and2 gate( .a(N2989), .b(EX677), .O(EX678) );
or2  gate( .a(EX672), .b(EX674), .O(EX679) );
or2  gate( .a(EX676), .b(EX679), .O(EX680) );
or2  gate( .a(EX678), .b(EX680), .O(N3212) );
and2 gate787( .a(N128), .b(N2990), .O(N3213) );
and2 gate788( .a(N125), .b(N2991), .O(N3214) );
and2 gate789( .a(N125), .b(N2992), .O(N3215) );
and2 gate790( .a(N655), .b(N2993), .O(N3216) );
inv1 gate( .a(N159),.O(N159_NOT) );
inv1 gate( .a(N2994),.O(N2994_NOT));
and2 gate( .a(N159_NOT), .b(p273), .O(EX681) );
and2 gate( .a(N2994_NOT), .b(EX681), .O(EX682) );
and2 gate( .a(N159), .b(p274), .O(EX683) );
and2 gate( .a(N2994_NOT), .b(EX683), .O(EX684) );
and2 gate( .a(N159_NOT), .b(p275), .O(EX685) );
and2 gate( .a(N2994), .b(EX685), .O(EX686) );
and2 gate( .a(N159), .b(p276), .O(EX687) );
and2 gate( .a(N2994), .b(EX687), .O(EX688) );
or2  gate( .a(EX682), .b(EX684), .O(EX689) );
or2  gate( .a(EX686), .b(EX689), .O(EX690) );
or2  gate( .a(EX688), .b(EX690), .O(N3217) );
and2 gate792( .a(N150), .b(N2995), .O(N3218) );
and2 gate793( .a(N143), .b(N2996), .O(N3219) );
and2 gate794( .a(N137), .b(N2997), .O(N3220) );
and2 gate795( .a(N132), .b(N2998), .O(N3221) );
and2 gate796( .a(N128), .b(N2999), .O(N3222) );
and2 gate797( .a(N128), .b(N3000), .O(N3223) );
and2 gate798( .a(N670), .b(N3001), .O(N3224) );
and2 gate799( .a(N655), .b(N3002), .O(N3225) );
and2 gate800( .a(N159), .b(N3003), .O(N3226) );
and2 gate801( .a(N150), .b(N3004), .O(N3227) );
and2 gate802( .a(N143), .b(N3005), .O(N3228) );
and2 gate803( .a(N137), .b(N3006), .O(N3229) );
and2 gate804( .a(N132), .b(N3007), .O(N3230) );
and2 gate805( .a(N132), .b(N3008), .O(N3231) );
and2 gate806( .a(N690), .b(N3009), .O(N3232) );
and2 gate807( .a(N670), .b(N3010), .O(N3233) );
and2 gate808( .a(N655), .b(N3011), .O(N3234) );
and2 gate809( .a(N159), .b(N3012), .O(N3235) );
and2 gate810( .a(N150), .b(N3013), .O(N3236) );
and2 gate811( .a(N143), .b(N3014), .O(N3237) );
and2 gate812( .a(N137), .b(N3015), .O(N3238) );
and2 gate813( .a(N137), .b(N3016), .O(N3239) );
and2 gate814( .a(N706), .b(N3017), .O(N3240) );
and2 gate815( .a(N690), .b(N3018), .O(N3241) );
and2 gate816( .a(N670), .b(N3019), .O(N3242) );
inv1 gate( .a(N655),.O(N655_NOT) );
inv1 gate( .a(N3020),.O(N3020_NOT));
and2 gate( .a(N655_NOT), .b(p277), .O(EX691) );
and2 gate( .a(N3020_NOT), .b(EX691), .O(EX692) );
and2 gate( .a(N655), .b(p278), .O(EX693) );
and2 gate( .a(N3020_NOT), .b(EX693), .O(EX694) );
and2 gate( .a(N655_NOT), .b(p279), .O(EX695) );
and2 gate( .a(N3020), .b(EX695), .O(EX696) );
and2 gate( .a(N655), .b(p280), .O(EX697) );
and2 gate( .a(N3020), .b(EX697), .O(EX698) );
or2  gate( .a(EX692), .b(EX694), .O(EX699) );
or2  gate( .a(EX696), .b(EX699), .O(EX700) );
or2  gate( .a(EX698), .b(EX700), .O(N3243) );
and2 gate818( .a(N159), .b(N3021), .O(N3244) );
and2 gate819( .a(N150), .b(N3022), .O(N3245) );
and2 gate820( .a(N143), .b(N3023), .O(N3246) );
and2 gate821( .a(N143), .b(N3024), .O(N3247) );
inv1 gate( .a(N715),.O(N715_NOT) );
inv1 gate( .a(N3025),.O(N3025_NOT));
and2 gate( .a(N715_NOT), .b(p281), .O(EX701) );
and2 gate( .a(N3025_NOT), .b(EX701), .O(EX702) );
and2 gate( .a(N715), .b(p282), .O(EX703) );
and2 gate( .a(N3025_NOT), .b(EX703), .O(EX704) );
and2 gate( .a(N715_NOT), .b(p283), .O(EX705) );
and2 gate( .a(N3025), .b(EX705), .O(EX706) );
and2 gate( .a(N715), .b(p284), .O(EX707) );
and2 gate( .a(N3025), .b(EX707), .O(EX708) );
or2  gate( .a(EX702), .b(EX704), .O(EX709) );
or2  gate( .a(EX706), .b(EX709), .O(EX710) );
or2  gate( .a(EX708), .b(EX710), .O(N3248) );
and2 gate823( .a(N706), .b(N3026), .O(N3249) );
and2 gate824( .a(N690), .b(N3027), .O(N3250) );
inv1 gate( .a(N670),.O(N670_NOT) );
inv1 gate( .a(N3028),.O(N3028_NOT));
and2 gate( .a(N670_NOT), .b(p285), .O(EX711) );
and2 gate( .a(N3028_NOT), .b(EX711), .O(EX712) );
and2 gate( .a(N670), .b(p286), .O(EX713) );
and2 gate( .a(N3028_NOT), .b(EX713), .O(EX714) );
and2 gate( .a(N670_NOT), .b(p287), .O(EX715) );
and2 gate( .a(N3028), .b(EX715), .O(EX716) );
and2 gate( .a(N670), .b(p288), .O(EX717) );
and2 gate( .a(N3028), .b(EX717), .O(EX718) );
or2  gate( .a(EX712), .b(EX714), .O(EX719) );
or2  gate( .a(EX716), .b(EX719), .O(EX720) );
or2  gate( .a(EX718), .b(EX720), .O(N3251) );
and2 gate826( .a(N655), .b(N3029), .O(N3252) );
and2 gate827( .a(N159), .b(N3030), .O(N3253) );
and2 gate828( .a(N150), .b(N3031), .O(N3254) );
inv1 gate( .a(N150),.O(N150_NOT) );
inv1 gate( .a(N3032),.O(N3032_NOT));
and2 gate( .a(N150_NOT), .b(p289), .O(EX721) );
and2 gate( .a(N3032_NOT), .b(EX721), .O(EX722) );
and2 gate( .a(N150), .b(p290), .O(EX723) );
and2 gate( .a(N3032_NOT), .b(EX723), .O(EX724) );
and2 gate( .a(N150_NOT), .b(p291), .O(EX725) );
and2 gate( .a(N3032), .b(EX725), .O(EX726) );
and2 gate( .a(N150), .b(p292), .O(EX727) );
and2 gate( .a(N3032), .b(EX727), .O(EX728) );
or2  gate( .a(EX722), .b(EX724), .O(EX729) );
or2  gate( .a(EX726), .b(EX729), .O(EX730) );
or2  gate( .a(EX728), .b(EX730), .O(N3255) );
and2 gate830( .a(N727), .b(N3033), .O(N3256) );
and2 gate831( .a(N715), .b(N3034), .O(N3257) );
and2 gate832( .a(N706), .b(N3035), .O(N3258) );
inv1 gate( .a(N690),.O(N690_NOT) );
inv1 gate( .a(N3036),.O(N3036_NOT));
and2 gate( .a(N690_NOT), .b(p293), .O(EX731) );
and2 gate( .a(N3036_NOT), .b(EX731), .O(EX732) );
and2 gate( .a(N690), .b(p294), .O(EX733) );
and2 gate( .a(N3036_NOT), .b(EX733), .O(EX734) );
and2 gate( .a(N690_NOT), .b(p295), .O(EX735) );
and2 gate( .a(N3036), .b(EX735), .O(EX736) );
and2 gate( .a(N690), .b(p296), .O(EX737) );
and2 gate( .a(N3036), .b(EX737), .O(EX738) );
or2  gate( .a(EX732), .b(EX734), .O(EX739) );
or2  gate( .a(EX736), .b(EX739), .O(EX740) );
or2  gate( .a(EX738), .b(EX740), .O(N3259) );
and2 gate834( .a(N670), .b(N3037), .O(N3260) );
and2 gate835( .a(N655), .b(N3038), .O(N3261) );
and2 gate836( .a(N159), .b(N3039), .O(N3262) );
and2 gate837( .a(N159), .b(N3040), .O(N3263) );
and2 gate838( .a(N740), .b(N3041), .O(N3264) );
and2 gate839( .a(N727), .b(N3042), .O(N3265) );
and2 gate840( .a(N715), .b(N3043), .O(N3266) );
and2 gate841( .a(N706), .b(N3044), .O(N3267) );
and2 gate842( .a(N690), .b(N3045), .O(N3268) );
and2 gate843( .a(N670), .b(N3046), .O(N3269) );
and2 gate844( .a(N655), .b(N3047), .O(N3270) );
inv1 gate( .a(N283),.O(N283_NOT) );
inv1 gate( .a(N3048),.O(N3048_NOT));
and2 gate( .a(N283_NOT), .b(p297), .O(EX741) );
and2 gate( .a(N3048_NOT), .b(EX741), .O(EX742) );
and2 gate( .a(N283), .b(p298), .O(EX743) );
and2 gate( .a(N3048_NOT), .b(EX743), .O(EX744) );
and2 gate( .a(N283_NOT), .b(p299), .O(EX745) );
and2 gate( .a(N3048), .b(EX745), .O(EX746) );
and2 gate( .a(N283), .b(p300), .O(EX747) );
and2 gate( .a(N3048), .b(EX747), .O(EX748) );
or2  gate( .a(EX742), .b(EX744), .O(EX749) );
or2  gate( .a(EX746), .b(EX749), .O(EX750) );
or2  gate( .a(EX748), .b(EX750), .O(N3271) );
and2 gate846( .a(N670), .b(N3049), .O(N3272) );
and2 gate847( .a(N690), .b(N3050), .O(N3273) );
and2 gate848( .a(N706), .b(N3051), .O(N3274) );
and2 gate849( .a(N715), .b(N3052), .O(N3275) );
inv1 gate( .a(N727),.O(N727_NOT) );
inv1 gate( .a(N3053),.O(N3053_NOT));
and2 gate( .a(N727_NOT), .b(p301), .O(EX751) );
and2 gate( .a(N3053_NOT), .b(EX751), .O(EX752) );
and2 gate( .a(N727), .b(p302), .O(EX753) );
and2 gate( .a(N3053_NOT), .b(EX753), .O(EX754) );
and2 gate( .a(N727_NOT), .b(p303), .O(EX755) );
and2 gate( .a(N3053), .b(EX755), .O(EX756) );
and2 gate( .a(N727), .b(p304), .O(EX757) );
and2 gate( .a(N3053), .b(EX757), .O(EX758) );
or2  gate( .a(EX752), .b(EX754), .O(EX759) );
or2  gate( .a(EX756), .b(EX759), .O(EX760) );
or2  gate( .a(EX758), .b(EX760), .O(N3276) );
and2 gate851( .a(N740), .b(N3054), .O(N3277) );
and2 gate852( .a(N753), .b(N3055), .O(N3278) );
and2 gate853( .a(N294), .b(N3056), .O(N3279) );
and2 gate854( .a(N690), .b(N3057), .O(N3280) );
and2 gate855( .a(N706), .b(N3058), .O(N3281) );
and2 gate856( .a(N715), .b(N3059), .O(N3282) );
and2 gate857( .a(N727), .b(N3060), .O(N3283) );
and2 gate858( .a(N740), .b(N3061), .O(N3284) );
inv1 gate( .a(N753),.O(N753_NOT) );
inv1 gate( .a(N3062),.O(N3062_NOT));
and2 gate( .a(N753_NOT), .b(p305), .O(EX761) );
and2 gate( .a(N3062_NOT), .b(EX761), .O(EX762) );
and2 gate( .a(N753), .b(p306), .O(EX763) );
and2 gate( .a(N3062_NOT), .b(EX763), .O(EX764) );
and2 gate( .a(N753_NOT), .b(p307), .O(EX765) );
and2 gate( .a(N3062), .b(EX765), .O(EX766) );
and2 gate( .a(N753), .b(p308), .O(EX767) );
and2 gate( .a(N3062), .b(EX767), .O(EX768) );
or2  gate( .a(EX762), .b(EX764), .O(EX769) );
or2  gate( .a(EX766), .b(EX769), .O(EX770) );
or2  gate( .a(EX768), .b(EX770), .O(N3285) );
inv1 gate( .a(N283),.O(N283_NOT) );
inv1 gate( .a(N3063),.O(N3063_NOT));
and2 gate( .a(N283_NOT), .b(p309), .O(EX771) );
and2 gate( .a(N3063_NOT), .b(EX771), .O(EX772) );
and2 gate( .a(N283), .b(p310), .O(EX773) );
and2 gate( .a(N3063_NOT), .b(EX773), .O(EX774) );
and2 gate( .a(N283_NOT), .b(p311), .O(EX775) );
and2 gate( .a(N3063), .b(EX775), .O(EX776) );
and2 gate( .a(N283), .b(p312), .O(EX777) );
and2 gate( .a(N3063), .b(EX777), .O(EX778) );
or2  gate( .a(EX772), .b(EX774), .O(EX779) );
or2  gate( .a(EX776), .b(EX779), .O(EX780) );
or2  gate( .a(EX778), .b(EX780), .O(N3286) );
and2 gate861( .a(N303), .b(N3064), .O(N3287) );
and2 gate862( .a(N706), .b(N3065), .O(N3288) );
inv1 gate( .a(N715),.O(N715_NOT) );
inv1 gate( .a(N3066),.O(N3066_NOT));
and2 gate( .a(N715_NOT), .b(p313), .O(EX781) );
and2 gate( .a(N3066_NOT), .b(EX781), .O(EX782) );
and2 gate( .a(N715), .b(p314), .O(EX783) );
and2 gate( .a(N3066_NOT), .b(EX783), .O(EX784) );
and2 gate( .a(N715_NOT), .b(p315), .O(EX785) );
and2 gate( .a(N3066), .b(EX785), .O(EX786) );
and2 gate( .a(N715), .b(p316), .O(EX787) );
and2 gate( .a(N3066), .b(EX787), .O(EX788) );
or2  gate( .a(EX782), .b(EX784), .O(EX789) );
or2  gate( .a(EX786), .b(EX789), .O(EX790) );
or2  gate( .a(EX788), .b(EX790), .O(N3289) );
and2 gate864( .a(N727), .b(N3067), .O(N3290) );
inv1 gate( .a(N740),.O(N740_NOT) );
inv1 gate( .a(N3068),.O(N3068_NOT));
and2 gate( .a(N740_NOT), .b(p317), .O(EX791) );
and2 gate( .a(N3068_NOT), .b(EX791), .O(EX792) );
and2 gate( .a(N740), .b(p318), .O(EX793) );
and2 gate( .a(N3068_NOT), .b(EX793), .O(EX794) );
and2 gate( .a(N740_NOT), .b(p319), .O(EX795) );
and2 gate( .a(N3068), .b(EX795), .O(EX796) );
and2 gate( .a(N740), .b(p320), .O(EX797) );
and2 gate( .a(N3068), .b(EX797), .O(EX798) );
or2  gate( .a(EX792), .b(EX794), .O(EX799) );
or2  gate( .a(EX796), .b(EX799), .O(EX800) );
or2  gate( .a(EX798), .b(EX800), .O(N3291) );
and2 gate866( .a(N753), .b(N3069), .O(N3292) );
and2 gate867( .a(N283), .b(N3070), .O(N3293) );
and2 gate868( .a(N294), .b(N3071), .O(N3294) );
inv1 gate( .a(N311),.O(N311_NOT) );
inv1 gate( .a(N3072),.O(N3072_NOT));
and2 gate( .a(N311_NOT), .b(p321), .O(EX801) );
and2 gate( .a(N3072_NOT), .b(EX801), .O(EX802) );
and2 gate( .a(N311), .b(p322), .O(EX803) );
and2 gate( .a(N3072_NOT), .b(EX803), .O(EX804) );
and2 gate( .a(N311_NOT), .b(p323), .O(EX805) );
and2 gate( .a(N3072), .b(EX805), .O(EX806) );
and2 gate( .a(N311), .b(p324), .O(EX807) );
and2 gate( .a(N3072), .b(EX807), .O(EX808) );
or2  gate( .a(EX802), .b(EX804), .O(EX809) );
or2  gate( .a(EX806), .b(EX809), .O(EX810) );
or2  gate( .a(EX808), .b(EX810), .O(N3295) );
inv1 gate( .a(N715),.O(N715_NOT) );
inv1 gate( .a(N3073),.O(N3073_NOT));
and2 gate( .a(N715_NOT), .b(p325), .O(EX811) );
and2 gate( .a(N3073_NOT), .b(EX811), .O(EX812) );
and2 gate( .a(N715), .b(p326), .O(EX813) );
and2 gate( .a(N3073_NOT), .b(EX813), .O(EX814) );
and2 gate( .a(N715_NOT), .b(p327), .O(EX815) );
and2 gate( .a(N3073), .b(EX815), .O(EX816) );
and2 gate( .a(N715), .b(p328), .O(EX817) );
and2 gate( .a(N3073), .b(EX817), .O(EX818) );
or2  gate( .a(EX812), .b(EX814), .O(EX819) );
or2  gate( .a(EX816), .b(EX819), .O(EX820) );
or2  gate( .a(EX818), .b(EX820), .O(N3296) );
inv1 gate( .a(N727),.O(N727_NOT) );
inv1 gate( .a(N3074),.O(N3074_NOT));
and2 gate( .a(N727_NOT), .b(p329), .O(EX821) );
and2 gate( .a(N3074_NOT), .b(EX821), .O(EX822) );
and2 gate( .a(N727), .b(p330), .O(EX823) );
and2 gate( .a(N3074_NOT), .b(EX823), .O(EX824) );
and2 gate( .a(N727_NOT), .b(p331), .O(EX825) );
and2 gate( .a(N3074), .b(EX825), .O(EX826) );
and2 gate( .a(N727), .b(p332), .O(EX827) );
and2 gate( .a(N3074), .b(EX827), .O(EX828) );
or2  gate( .a(EX822), .b(EX824), .O(EX829) );
or2  gate( .a(EX826), .b(EX829), .O(EX830) );
or2  gate( .a(EX828), .b(EX830), .O(N3297) );
inv1 gate( .a(N740),.O(N740_NOT) );
inv1 gate( .a(N3075),.O(N3075_NOT));
and2 gate( .a(N740_NOT), .b(p333), .O(EX831) );
and2 gate( .a(N3075_NOT), .b(EX831), .O(EX832) );
and2 gate( .a(N740), .b(p334), .O(EX833) );
and2 gate( .a(N3075_NOT), .b(EX833), .O(EX834) );
and2 gate( .a(N740_NOT), .b(p335), .O(EX835) );
and2 gate( .a(N3075), .b(EX835), .O(EX836) );
and2 gate( .a(N740), .b(p336), .O(EX837) );
and2 gate( .a(N3075), .b(EX837), .O(EX838) );
or2  gate( .a(EX832), .b(EX834), .O(EX839) );
or2  gate( .a(EX836), .b(EX839), .O(EX840) );
or2  gate( .a(EX838), .b(EX840), .O(N3298) );
and2 gate873( .a(N753), .b(N3076), .O(N3299) );
and2 gate874( .a(N283), .b(N3077), .O(N3300) );
and2 gate875( .a(N294), .b(N3078), .O(N3301) );
and2 gate876( .a(N303), .b(N3079), .O(N3302) );
inv1 gate( .a(N317),.O(N317_NOT) );
inv1 gate( .a(N3080),.O(N3080_NOT));
and2 gate( .a(N317_NOT), .b(p337), .O(EX841) );
and2 gate( .a(N3080_NOT), .b(EX841), .O(EX842) );
and2 gate( .a(N317), .b(p338), .O(EX843) );
and2 gate( .a(N3080_NOT), .b(EX843), .O(EX844) );
and2 gate( .a(N317_NOT), .b(p339), .O(EX845) );
and2 gate( .a(N3080), .b(EX845), .O(EX846) );
and2 gate( .a(N317), .b(p340), .O(EX847) );
and2 gate( .a(N3080), .b(EX847), .O(EX848) );
or2  gate( .a(EX842), .b(EX844), .O(EX849) );
or2  gate( .a(EX846), .b(EX849), .O(EX850) );
or2  gate( .a(EX848), .b(EX850), .O(N3303) );
and2 gate878( .a(N727), .b(N3081), .O(N3304) );
and2 gate879( .a(N740), .b(N3082), .O(N3305) );
and2 gate880( .a(N753), .b(N3083), .O(N3306) );
inv1 gate( .a(N283),.O(N283_NOT) );
inv1 gate( .a(N3084),.O(N3084_NOT));
and2 gate( .a(N283_NOT), .b(p341), .O(EX851) );
and2 gate( .a(N3084_NOT), .b(EX851), .O(EX852) );
and2 gate( .a(N283), .b(p342), .O(EX853) );
and2 gate( .a(N3084_NOT), .b(EX853), .O(EX854) );
and2 gate( .a(N283_NOT), .b(p343), .O(EX855) );
and2 gate( .a(N3084), .b(EX855), .O(EX856) );
and2 gate( .a(N283), .b(p344), .O(EX857) );
and2 gate( .a(N3084), .b(EX857), .O(EX858) );
or2  gate( .a(EX852), .b(EX854), .O(EX859) );
or2  gate( .a(EX856), .b(EX859), .O(EX860) );
or2  gate( .a(EX858), .b(EX860), .O(N3307) );
inv1 gate( .a(N294),.O(N294_NOT) );
inv1 gate( .a(N3085),.O(N3085_NOT));
and2 gate( .a(N294_NOT), .b(p345), .O(EX861) );
and2 gate( .a(N3085_NOT), .b(EX861), .O(EX862) );
and2 gate( .a(N294), .b(p346), .O(EX863) );
and2 gate( .a(N3085_NOT), .b(EX863), .O(EX864) );
and2 gate( .a(N294_NOT), .b(p347), .O(EX865) );
and2 gate( .a(N3085), .b(EX865), .O(EX866) );
and2 gate( .a(N294), .b(p348), .O(EX867) );
and2 gate( .a(N3085), .b(EX867), .O(EX868) );
or2  gate( .a(EX862), .b(EX864), .O(EX869) );
or2  gate( .a(EX866), .b(EX869), .O(EX870) );
or2  gate( .a(EX868), .b(EX870), .O(N3308) );
and2 gate883( .a(N303), .b(N3086), .O(N3309) );
and2 gate884( .a(N311), .b(N3087), .O(N3310) );
and2 gate885( .a(N322), .b(N3088), .O(N3311) );
and2 gate886( .a(N740), .b(N3089), .O(N3312) );
inv1 gate( .a(N753),.O(N753_NOT) );
inv1 gate( .a(N3090),.O(N3090_NOT));
and2 gate( .a(N753_NOT), .b(p349), .O(EX871) );
and2 gate( .a(N3090_NOT), .b(EX871), .O(EX872) );
and2 gate( .a(N753), .b(p350), .O(EX873) );
and2 gate( .a(N3090_NOT), .b(EX873), .O(EX874) );
and2 gate( .a(N753_NOT), .b(p351), .O(EX875) );
and2 gate( .a(N3090), .b(EX875), .O(EX876) );
and2 gate( .a(N753), .b(p352), .O(EX877) );
and2 gate( .a(N3090), .b(EX877), .O(EX878) );
or2  gate( .a(EX872), .b(EX874), .O(EX879) );
or2  gate( .a(EX876), .b(EX879), .O(EX880) );
or2  gate( .a(EX878), .b(EX880), .O(N3313) );
inv1 gate( .a(N283),.O(N283_NOT) );
inv1 gate( .a(N3091),.O(N3091_NOT));
and2 gate( .a(N283_NOT), .b(p353), .O(EX881) );
and2 gate( .a(N3091_NOT), .b(EX881), .O(EX882) );
and2 gate( .a(N283), .b(p354), .O(EX883) );
and2 gate( .a(N3091_NOT), .b(EX883), .O(EX884) );
and2 gate( .a(N283_NOT), .b(p355), .O(EX885) );
and2 gate( .a(N3091), .b(EX885), .O(EX886) );
and2 gate( .a(N283), .b(p356), .O(EX887) );
and2 gate( .a(N3091), .b(EX887), .O(EX888) );
or2  gate( .a(EX882), .b(EX884), .O(EX889) );
or2  gate( .a(EX886), .b(EX889), .O(EX890) );
or2  gate( .a(EX888), .b(EX890), .O(N3314) );
and2 gate889( .a(N294), .b(N3092), .O(N3315) );
inv1 gate( .a(N303),.O(N303_NOT) );
inv1 gate( .a(N3093),.O(N3093_NOT));
and2 gate( .a(N303_NOT), .b(p357), .O(EX891) );
and2 gate( .a(N3093_NOT), .b(EX891), .O(EX892) );
and2 gate( .a(N303), .b(p358), .O(EX893) );
and2 gate( .a(N3093_NOT), .b(EX893), .O(EX894) );
and2 gate( .a(N303_NOT), .b(p359), .O(EX895) );
and2 gate( .a(N3093), .b(EX895), .O(EX896) );
and2 gate( .a(N303), .b(p360), .O(EX897) );
and2 gate( .a(N3093), .b(EX897), .O(EX898) );
or2  gate( .a(EX892), .b(EX894), .O(EX899) );
or2  gate( .a(EX896), .b(EX899), .O(EX900) );
or2  gate( .a(EX898), .b(EX900), .O(N3316) );
and2 gate891( .a(N311), .b(N3094), .O(N3317) );
inv1 gate( .a(N317),.O(N317_NOT) );
inv1 gate( .a(N3095),.O(N3095_NOT));
and2 gate( .a(N317_NOT), .b(p361), .O(EX901) );
and2 gate( .a(N3095_NOT), .b(EX901), .O(EX902) );
and2 gate( .a(N317), .b(p362), .O(EX903) );
and2 gate( .a(N3095_NOT), .b(EX903), .O(EX904) );
and2 gate( .a(N317_NOT), .b(p363), .O(EX905) );
and2 gate( .a(N3095), .b(EX905), .O(EX906) );
and2 gate( .a(N317), .b(p364), .O(EX907) );
and2 gate( .a(N3095), .b(EX907), .O(EX908) );
or2  gate( .a(EX902), .b(EX904), .O(EX909) );
or2  gate( .a(EX906), .b(EX909), .O(EX910) );
or2  gate( .a(EX908), .b(EX910), .O(N3318) );
and2 gate893( .a(N326), .b(N3096), .O(N3319) );
and2 gate894( .a(N753), .b(N3097), .O(N3320) );
inv1 gate( .a(N283),.O(N283_NOT) );
inv1 gate( .a(N3098),.O(N3098_NOT));
and2 gate( .a(N283_NOT), .b(p365), .O(EX911) );
and2 gate( .a(N3098_NOT), .b(EX911), .O(EX912) );
and2 gate( .a(N283), .b(p366), .O(EX913) );
and2 gate( .a(N3098_NOT), .b(EX913), .O(EX914) );
and2 gate( .a(N283_NOT), .b(p367), .O(EX915) );
and2 gate( .a(N3098), .b(EX915), .O(EX916) );
and2 gate( .a(N283), .b(p368), .O(EX917) );
and2 gate( .a(N3098), .b(EX917), .O(EX918) );
or2  gate( .a(EX912), .b(EX914), .O(EX919) );
or2  gate( .a(EX916), .b(EX919), .O(EX920) );
or2  gate( .a(EX918), .b(EX920), .O(N3321) );
and2 gate896( .a(N294), .b(N3099), .O(N3322) );
and2 gate897( .a(N303), .b(N3100), .O(N3323) );
and2 gate898( .a(N311), .b(N3101), .O(N3324) );
and2 gate899( .a(N317), .b(N3102), .O(N3325) );
and2 gate900( .a(N322), .b(N3103), .O(N3326) );
inv1 gate( .a(N329),.O(N329_NOT) );
inv1 gate( .a(N3104),.O(N3104_NOT));
and2 gate( .a(N329_NOT), .b(p369), .O(EX921) );
and2 gate( .a(N3104_NOT), .b(EX921), .O(EX922) );
and2 gate( .a(N329), .b(p370), .O(EX923) );
and2 gate( .a(N3104_NOT), .b(EX923), .O(EX924) );
and2 gate( .a(N329_NOT), .b(p371), .O(EX925) );
and2 gate( .a(N3104), .b(EX925), .O(EX926) );
and2 gate( .a(N329), .b(p372), .O(EX927) );
and2 gate( .a(N3104), .b(EX927), .O(EX928) );
or2  gate( .a(EX922), .b(EX924), .O(EX929) );
or2  gate( .a(EX926), .b(EX929), .O(EX930) );
or2  gate( .a(EX928), .b(EX930), .O(N3327) );
and2 gate902( .a(N283), .b(N3105), .O(N3328) );
and2 gate903( .a(N294), .b(N3106), .O(N3329) );
and2 gate904( .a(N303), .b(N3107), .O(N3330) );
and2 gate905( .a(N311), .b(N3108), .O(N3331) );
and2 gate906( .a(N317), .b(N3109), .O(N3332) );
and2 gate907( .a(N322), .b(N3110), .O(N3333) );
and2 gate908( .a(N326), .b(N3111), .O(N3334) );
and5 gate909( .a(N3190), .b(N3191), .c(N3192), .d(N3193), .e(N917), .O(N3383) );
buf1 gate910( .a(N2977), .O(N3384) );
inv1 gate( .a(N3196),.O(N3196_NOT) );
inv1 gate( .a(N1736),.O(N1736_NOT));
and2 gate( .a(N3196_NOT), .b(p373), .O(EX931) );
and2 gate( .a(N1736_NOT), .b(EX931), .O(EX932) );
and2 gate( .a(N3196), .b(p374), .O(EX933) );
and2 gate( .a(N1736_NOT), .b(EX933), .O(EX934) );
and2 gate( .a(N3196_NOT), .b(p375), .O(EX935) );
and2 gate( .a(N1736), .b(EX935), .O(EX936) );
and2 gate( .a(N3196), .b(p376), .O(EX937) );
and2 gate( .a(N1736), .b(EX937), .O(EX938) );
or2  gate( .a(EX932), .b(EX934), .O(EX939) );
or2  gate( .a(EX936), .b(EX939), .O(EX940) );
or2  gate( .a(EX938), .b(EX940), .O(N3387) );
and2 gate912( .a(N2977), .b(N2149), .O(N3388) );
and2 gate913( .a(N2973), .b(N1737), .O(N3389) );
nor8 gate914( .a(N3207), .b(N3208), .c(N3209), .d(N3210), .e(N3211), .f(N3212), .g(N3213), .h(N3214), .O(N3390) );
nor8 gate915( .a(N3215), .b(N3216), .c(N3217), .d(N3218), .e(N3219), .f(N3220), .g(N3221), .h(N3222), .O(N3391) );
nor8 gate916( .a(N3223), .b(N3224), .c(N3225), .d(N3226), .e(N3227), .f(N3228), .g(N3229), .h(N3230), .O(N3392) );
nor8 gate917( .a(N3231), .b(N3232), .c(N3233), .d(N3234), .e(N3235), .f(N3236), .g(N3237), .h(N3238), .O(N3393) );
nor8 gate918( .a(N3239), .b(N3240), .c(N3241), .d(N3242), .e(N3243), .f(N3244), .g(N3245), .h(N3246), .O(N3394) );
nor8 gate919( .a(N3247), .b(N3248), .c(N3249), .d(N3250), .e(N3251), .f(N3252), .g(N3253), .h(N3254), .O(N3395) );
nor8 gate920( .a(N3255), .b(N3256), .c(N3257), .d(N3258), .e(N3259), .f(N3260), .g(N3261), .h(N3262), .O(N3396) );
nor8 gate921( .a(N3263), .b(N3264), .c(N3265), .d(N3266), .e(N3267), .f(N3268), .g(N3269), .h(N3270), .O(N3397) );
nor8 gate922( .a(N3271), .b(N3272), .c(N3273), .d(N3274), .e(N3275), .f(N3276), .g(N3277), .h(N3278), .O(N3398) );
nor8 gate923( .a(N3279), .b(N3280), .c(N3281), .d(N3282), .e(N3283), .f(N3284), .g(N3285), .h(N3286), .O(N3399) );
nor8 gate924( .a(N3287), .b(N3288), .c(N3289), .d(N3290), .e(N3291), .f(N3292), .g(N3293), .h(N3294), .O(N3400) );
nor8 gate925( .a(N3295), .b(N3296), .c(N3297), .d(N3298), .e(N3299), .f(N3300), .g(N3301), .h(N3302), .O(N3401) );
nor8 gate926( .a(N3303), .b(N3304), .c(N3305), .d(N3306), .e(N3307), .f(N3308), .g(N3309), .h(N3310), .O(N3402) );
nor8 gate927( .a(N3311), .b(N3312), .c(N3313), .d(N3314), .e(N3315), .f(N3316), .g(N3317), .h(N3318), .O(N3403) );
nor8 gate928( .a(N3319), .b(N3320), .c(N3321), .d(N3322), .e(N3323), .f(N3324), .g(N3325), .h(N3326), .O(N3404) );
nor8 gate929( .a(N3327), .b(N3328), .c(N3329), .d(N3330), .e(N3331), .f(N3332), .g(N3333), .h(N3334), .O(N3405) );
and2 gate930( .a(N3206), .b(N2641), .O(N3406) );
and3 gate931( .a(N169), .b(N2648), .c(N3112), .O(N3407) );
and3 gate932( .a(N179), .b(N2648), .c(N3115), .O(N3410) );
and3 gate933( .a(N190), .b(N2652), .c(N3115), .O(N3413) );
and3 gate934( .a(N200), .b(N2652), .c(N3112), .O(N3414) );
or3 gate935( .a(N3119), .b(N1875), .c(N2073), .O(N3415) );
nor3 gate936( .a(N3119), .b(N1875), .c(N2073), .O(N3419) );
and3 gate937( .a(N169), .b(N2662), .c(N3128), .O(N3423) );
and3 gate938( .a(N179), .b(N2662), .c(N3131), .O(N3426) );
and3 gate939( .a(N190), .b(N2666), .c(N3131), .O(N3429) );
and3 gate940( .a(N200), .b(N2666), .c(N3128), .O(N3430) );
and3 gate941( .a(N169), .b(N2673), .c(N3135), .O(N3431) );
and3 gate942( .a(N179), .b(N2673), .c(N3138), .O(N3434) );
and3 gate943( .a(N190), .b(N2677), .c(N3138), .O(N3437) );
and3 gate944( .a(N200), .b(N2677), .c(N3135), .O(N3438) );
and3 gate945( .a(N169), .b(N2684), .c(N3142), .O(N3439) );
and3 gate946( .a(N179), .b(N2684), .c(N3145), .O(N3442) );
and3 gate947( .a(N190), .b(N2688), .c(N3145), .O(N3445) );
and3 gate948( .a(N200), .b(N2688), .c(N3142), .O(N3446) );
or3 gate949( .a(N3149), .b(N1895), .c(N2093), .O(N3447) );
nor3 gate950( .a(N3149), .b(N1895), .c(N2093), .O(N3451) );
and3 gate951( .a(N169), .b(N2702), .c(N3158), .O(N3455) );
and3 gate952( .a(N179), .b(N2702), .c(N3161), .O(N3458) );
and3 gate953( .a(N190), .b(N2706), .c(N3161), .O(N3461) );
and3 gate954( .a(N200), .b(N2706), .c(N3158), .O(N3462) );
and3 gate955( .a(N169), .b(N2715), .c(N3165), .O(N3463) );
and3 gate956( .a(N179), .b(N2715), .c(N3168), .O(N3466) );
and3 gate957( .a(N190), .b(N2719), .c(N3168), .O(N3469) );
and3 gate958( .a(N200), .b(N2719), .c(N3165), .O(N3470) );
or2 gate959( .a(N3194), .b(N3383), .O(N3471) );
buf1 gate960( .a(N2967), .O(N3472) );
buf1 gate961( .a(N2970), .O(N3475) );
buf1 gate962( .a(N2967), .O(N3478) );
buf1 gate963( .a(N2970), .O(N3481) );
buf1 gate964( .a(N2973), .O(N3484) );
buf1 gate965( .a(N2973), .O(N3487) );
buf1 gate966( .a(N3172), .O(N3490) );
buf1 gate967( .a(N3172), .O(N3493) );
buf1 gate968( .a(N3175), .O(N3496) );
buf1 gate969( .a(N3175), .O(N3499) );
buf1 gate970( .a(N3178), .O(N3502) );
buf1 gate971( .a(N3178), .O(N3505) );
buf1 gate972( .a(N3181), .O(N3508) );
buf1 gate973( .a(N3181), .O(N3511) );
buf1 gate974( .a(N3184), .O(N3514) );
buf1 gate975( .a(N3184), .O(N3517) );
buf1 gate976( .a(N3187), .O(N3520) );
buf1 gate977( .a(N3187), .O(N3523) );
inv1 gate( .a(N3387),.O(N3387_NOT) );
inv1 gate( .a(N2350),.O(N2350_NOT));
and2 gate( .a(N3387_NOT), .b(p377), .O(EX941) );
and2 gate( .a(N2350_NOT), .b(EX941), .O(EX942) );
and2 gate( .a(N3387), .b(p378), .O(EX943) );
and2 gate( .a(N2350_NOT), .b(EX943), .O(EX944) );
and2 gate( .a(N3387_NOT), .b(p379), .O(EX945) );
and2 gate( .a(N2350), .b(EX945), .O(EX946) );
and2 gate( .a(N3387), .b(p380), .O(EX947) );
and2 gate( .a(N2350), .b(EX947), .O(EX948) );
or2  gate( .a(EX942), .b(EX944), .O(EX949) );
or2  gate( .a(EX946), .b(EX949), .O(EX950) );
or2  gate( .a(EX948), .b(EX950), .O(N3534) );
or3 gate979( .a(N3388), .b(N2151), .c(N2351), .O(N3535) );
nor2 gate980( .a(N3389), .b(N1966), .O(N3536) );
and2 gate981( .a(N3390), .b(N2209), .O(N3537) );
and2 gate982( .a(N3398), .b(N2210), .O(N3538) );
and2 gate983( .a(N3391), .b(N1842), .O(N3539) );
and2 gate984( .a(N3399), .b(N1369), .O(N3540) );
inv1 gate( .a(N3392),.O(N3392_NOT) );
inv1 gate( .a(N1843),.O(N1843_NOT));
and2 gate( .a(N3392_NOT), .b(p381), .O(EX951) );
and2 gate( .a(N1843_NOT), .b(EX951), .O(EX952) );
and2 gate( .a(N3392), .b(p382), .O(EX953) );
and2 gate( .a(N1843_NOT), .b(EX953), .O(EX954) );
and2 gate( .a(N3392_NOT), .b(p383), .O(EX955) );
and2 gate( .a(N1843), .b(EX955), .O(EX956) );
and2 gate( .a(N3392), .b(p384), .O(EX957) );
and2 gate( .a(N1843), .b(EX957), .O(EX958) );
or2  gate( .a(EX952), .b(EX954), .O(EX959) );
or2  gate( .a(EX956), .b(EX959), .O(EX960) );
or2  gate( .a(EX958), .b(EX960), .O(N3541) );
and2 gate986( .a(N3400), .b(N1369), .O(N3542) );
and2 gate987( .a(N3393), .b(N1844), .O(N3543) );
and2 gate988( .a(N3401), .b(N1369), .O(N3544) );
and2 gate989( .a(N3394), .b(N1845), .O(N3545) );
and2 gate990( .a(N3402), .b(N1369), .O(N3546) );
and2 gate991( .a(N3395), .b(N1846), .O(N3547) );
and2 gate992( .a(N3403), .b(N1369), .O(N3548) );
inv1 gate( .a(N3396),.O(N3396_NOT) );
inv1 gate( .a(N1847),.O(N1847_NOT));
and2 gate( .a(N3396_NOT), .b(p385), .O(EX961) );
and2 gate( .a(N1847_NOT), .b(EX961), .O(EX962) );
and2 gate( .a(N3396), .b(p386), .O(EX963) );
and2 gate( .a(N1847_NOT), .b(EX963), .O(EX964) );
and2 gate( .a(N3396_NOT), .b(p387), .O(EX965) );
and2 gate( .a(N1847), .b(EX965), .O(EX966) );
and2 gate( .a(N3396), .b(p388), .O(EX967) );
and2 gate( .a(N1847), .b(EX967), .O(EX968) );
or2  gate( .a(EX962), .b(EX964), .O(EX969) );
or2  gate( .a(EX966), .b(EX969), .O(EX970) );
or2  gate( .a(EX968), .b(EX970), .O(N3549) );
and2 gate994( .a(N3404), .b(N1369), .O(N3550) );
and2 gate995( .a(N3397), .b(N1848), .O(N3551) );
and2 gate996( .a(N3405), .b(N1369), .O(N3552) );
or3 gate997( .a(N3413), .b(N3414), .c(N3118), .O(N3557) );
or3 gate998( .a(N3429), .b(N3430), .c(N3134), .O(N3568) );
or3 gate999( .a(N3437), .b(N3438), .c(N3141), .O(N3573) );
or3 gate1000( .a(N3445), .b(N3446), .c(N3148), .O(N3578) );
or3 gate1001( .a(N3461), .b(N3462), .c(N3164), .O(N3589) );
or3 gate1002( .a(N3469), .b(N3470), .c(N3171), .O(N3594) );
and2 gate1003( .a(N3471), .b(N2728), .O(N3605) );
inv1 gate1004( .a(N3478), .O(N3626) );
inv1 gate1005( .a(N3481), .O(N3627) );
inv1 gate1006( .a(N3487), .O(N3628) );
inv1 gate1007( .a(N3484), .O(N3629) );
inv1 gate1008( .a(N3472), .O(N3630) );
inv1 gate1009( .a(N3475), .O(N3631) );
and2 gate1010( .a(N3536), .b(N2152), .O(N3632) );
and2 gate1011( .a(N3534), .b(N2155), .O(N3633) );
or3 gate1012( .a(N3537), .b(N3538), .c(N2398), .O(N3634) );
or2 gate1013( .a(N3539), .b(N3540), .O(N3635) );
or2 gate1014( .a(N3541), .b(N3542), .O(N3636) );
or2 gate1015( .a(N3543), .b(N3544), .O(N3637) );
or2 gate1016( .a(N3545), .b(N3546), .O(N3638) );
or2 gate1017( .a(N3547), .b(N3548), .O(N3639) );
or2 gate1018( .a(N3549), .b(N3550), .O(N3640) );
or2 gate1019( .a(N3551), .b(N3552), .O(N3641) );
and2 gate1020( .a(N3535), .b(N2643), .O(N3642) );
inv1 gate( .a(N3407),.O(N3407_NOT) );
inv1 gate( .a(N3410),.O(N3410_NOT));
and2 gate( .a(N3407_NOT), .b(p389), .O(EX971) );
and2 gate( .a(N3410_NOT), .b(EX971), .O(EX972) );
and2 gate( .a(N3407), .b(p390), .O(EX973) );
and2 gate( .a(N3410_NOT), .b(EX973), .O(EX974) );
and2 gate( .a(N3407_NOT), .b(p391), .O(EX975) );
and2 gate( .a(N3410), .b(EX975), .O(EX976) );
and2 gate( .a(N3407), .b(p392), .O(EX977) );
and2 gate( .a(N3410), .b(EX977), .O(EX978) );
or2  gate( .a(EX972), .b(EX974), .O(EX979) );
or2  gate( .a(EX976), .b(EX979), .O(EX980) );
or2  gate( .a(EX978), .b(EX980), .O(N3643) );
nor2 gate1022( .a(N3407), .b(N3410), .O(N3644) );
and3 gate1023( .a(N169), .b(N3415), .c(N3122), .O(N3645) );
and3 gate1024( .a(N179), .b(N3415), .c(N3125), .O(N3648) );
and3 gate1025( .a(N190), .b(N3419), .c(N3125), .O(N3651) );
and3 gate1026( .a(N200), .b(N3419), .c(N3122), .O(N3652) );
inv1 gate1027( .a(N3419), .O(N3653) );
or2 gate1028( .a(N3423), .b(N3426), .O(N3654) );
nor2 gate1029( .a(N3423), .b(N3426), .O(N3657) );
or2 gate1030( .a(N3431), .b(N3434), .O(N3658) );
nor2 gate1031( .a(N3431), .b(N3434), .O(N3661) );
or2 gate1032( .a(N3439), .b(N3442), .O(N3662) );
inv1 gate( .a(N3439),.O(N3439_NOT) );
inv1 gate( .a(N3442),.O(N3442_NOT));
and2 gate( .a(N3439_NOT), .b(p393), .O(EX981) );
and2 gate( .a(N3442_NOT), .b(EX981), .O(EX982) );
and2 gate( .a(N3439), .b(p394), .O(EX983) );
and2 gate( .a(N3442_NOT), .b(EX983), .O(EX984) );
and2 gate( .a(N3439_NOT), .b(p395), .O(EX985) );
and2 gate( .a(N3442), .b(EX985), .O(EX986) );
and2 gate( .a(N3439), .b(p396), .O(EX987) );
and2 gate( .a(N3442), .b(EX987), .O(EX988) );
or2  gate( .a(EX982), .b(EX984), .O(EX989) );
or2  gate( .a(EX986), .b(EX989), .O(EX990) );
or2  gate( .a(EX988), .b(EX990), .O(N3663) );
and3 gate1034( .a(N169), .b(N3447), .c(N3152), .O(N3664) );
and3 gate1035( .a(N179), .b(N3447), .c(N3155), .O(N3667) );
and3 gate1036( .a(N190), .b(N3451), .c(N3155), .O(N3670) );
and3 gate1037( .a(N200), .b(N3451), .c(N3152), .O(N3671) );
inv1 gate1038( .a(N3451), .O(N3672) );
or2 gate1039( .a(N3455), .b(N3458), .O(N3673) );
nor2 gate1040( .a(N3455), .b(N3458), .O(N3676) );
or2 gate1041( .a(N3463), .b(N3466), .O(N3677) );
nor2 gate1042( .a(N3463), .b(N3466), .O(N3680) );
inv1 gate1043( .a(N3493), .O(N3681) );
and2 gate1044( .a(N1909), .b(N3415), .O(N3682) );
inv1 gate1045( .a(N3496), .O(N3685) );
inv1 gate1046( .a(N3499), .O(N3686) );
inv1 gate1047( .a(N3502), .O(N3687) );
inv1 gate1048( .a(N3505), .O(N3688) );
inv1 gate1049( .a(N3511), .O(N3689) );
and2 gate1050( .a(N1922), .b(N3447), .O(N3690) );
inv1 gate1051( .a(N3517), .O(N3693) );
inv1 gate1052( .a(N3520), .O(N3694) );
inv1 gate1053( .a(N3523), .O(N3695) );
inv1 gate1054( .a(N3514), .O(N3696) );
buf1 gate1055( .a(N3384), .O(N3697) );
buf1 gate1056( .a(N3384), .O(N3700) );
inv1 gate1057( .a(N3490), .O(N3703) );
inv1 gate1058( .a(N3508), .O(N3704) );
inv1 gate( .a(N3475),.O(N3475_NOT) );
inv1 gate( .a(N3630),.O(N3630_NOT));
and2 gate( .a(N3475_NOT), .b(p397), .O(EX991) );
and2 gate( .a(N3630_NOT), .b(EX991), .O(EX992) );
and2 gate( .a(N3475), .b(p398), .O(EX993) );
and2 gate( .a(N3630_NOT), .b(EX993), .O(EX994) );
and2 gate( .a(N3475_NOT), .b(p399), .O(EX995) );
and2 gate( .a(N3630), .b(EX995), .O(EX996) );
and2 gate( .a(N3475), .b(p400), .O(EX997) );
and2 gate( .a(N3630), .b(EX997), .O(EX998) );
or2  gate( .a(EX992), .b(EX994), .O(EX999) );
or2  gate( .a(EX996), .b(EX999), .O(EX1000) );
or2  gate( .a(EX998), .b(EX1000), .O(N3705) );
nand2 gate1060( .a(N3472), .b(N3631), .O(N3706) );
inv1 gate( .a(N3481),.O(N3481_NOT) );
inv1 gate( .a(N3626),.O(N3626_NOT));
and2 gate( .a(N3481_NOT), .b(p401), .O(EX1001) );
and2 gate( .a(N3626_NOT), .b(EX1001), .O(EX1002) );
and2 gate( .a(N3481), .b(p402), .O(EX1003) );
and2 gate( .a(N3626_NOT), .b(EX1003), .O(EX1004) );
and2 gate( .a(N3481_NOT), .b(p403), .O(EX1005) );
and2 gate( .a(N3626), .b(EX1005), .O(EX1006) );
and2 gate( .a(N3481), .b(p404), .O(EX1007) );
and2 gate( .a(N3626), .b(EX1007), .O(EX1008) );
or2  gate( .a(EX1002), .b(EX1004), .O(EX1009) );
or2  gate( .a(EX1006), .b(EX1009), .O(EX1010) );
or2  gate( .a(EX1008), .b(EX1010), .O(N3707) );
inv1 gate( .a(N3478),.O(N3478_NOT) );
inv1 gate( .a(N3627),.O(N3627_NOT));
and2 gate( .a(N3478_NOT), .b(p405), .O(EX1011) );
and2 gate( .a(N3627_NOT), .b(EX1011), .O(EX1012) );
and2 gate( .a(N3478), .b(p406), .O(EX1013) );
and2 gate( .a(N3627_NOT), .b(EX1013), .O(EX1014) );
and2 gate( .a(N3478_NOT), .b(p407), .O(EX1015) );
and2 gate( .a(N3627), .b(EX1015), .O(EX1016) );
and2 gate( .a(N3478), .b(p408), .O(EX1017) );
and2 gate( .a(N3627), .b(EX1017), .O(EX1018) );
or2  gate( .a(EX1012), .b(EX1014), .O(EX1019) );
or2  gate( .a(EX1016), .b(EX1019), .O(EX1020) );
or2  gate( .a(EX1018), .b(EX1020), .O(N3708) );
or3 gate1063( .a(N3632), .b(N2352), .c(N2353), .O(N3711) );
or3 gate1064( .a(N3633), .b(N2354), .c(N2355), .O(N3712) );
and2 gate1065( .a(N3634), .b(N2632), .O(N3713) );
and2 gate1066( .a(N3635), .b(N2634), .O(N3714) );
inv1 gate( .a(N3636),.O(N3636_NOT) );
inv1 gate( .a(N2636),.O(N2636_NOT));
and2 gate( .a(N3636_NOT), .b(p409), .O(EX1021) );
and2 gate( .a(N2636_NOT), .b(EX1021), .O(EX1022) );
and2 gate( .a(N3636), .b(p410), .O(EX1023) );
and2 gate( .a(N2636_NOT), .b(EX1023), .O(EX1024) );
and2 gate( .a(N3636_NOT), .b(p411), .O(EX1025) );
and2 gate( .a(N2636), .b(EX1025), .O(EX1026) );
and2 gate( .a(N3636), .b(p412), .O(EX1027) );
and2 gate( .a(N2636), .b(EX1027), .O(EX1028) );
or2  gate( .a(EX1022), .b(EX1024), .O(EX1029) );
or2  gate( .a(EX1026), .b(EX1029), .O(EX1030) );
or2  gate( .a(EX1028), .b(EX1030), .O(N3715) );
inv1 gate( .a(N3637),.O(N3637_NOT) );
inv1 gate( .a(N2638),.O(N2638_NOT));
and2 gate( .a(N3637_NOT), .b(p413), .O(EX1031) );
and2 gate( .a(N2638_NOT), .b(EX1031), .O(EX1032) );
and2 gate( .a(N3637), .b(p414), .O(EX1033) );
and2 gate( .a(N2638_NOT), .b(EX1033), .O(EX1034) );
and2 gate( .a(N3637_NOT), .b(p415), .O(EX1035) );
and2 gate( .a(N2638), .b(EX1035), .O(EX1036) );
and2 gate( .a(N3637), .b(p416), .O(EX1037) );
and2 gate( .a(N2638), .b(EX1037), .O(EX1038) );
or2  gate( .a(EX1032), .b(EX1034), .O(EX1039) );
or2  gate( .a(EX1036), .b(EX1039), .O(EX1040) );
or2  gate( .a(EX1038), .b(EX1040), .O(N3716) );
and2 gate1069( .a(N3638), .b(N2640), .O(N3717) );
and2 gate1070( .a(N3639), .b(N2642), .O(N3718) );
and2 gate1071( .a(N3640), .b(N2644), .O(N3719) );
inv1 gate( .a(N3641),.O(N3641_NOT) );
inv1 gate( .a(N2646),.O(N2646_NOT));
and2 gate( .a(N3641_NOT), .b(p417), .O(EX1041) );
and2 gate( .a(N2646_NOT), .b(EX1041), .O(EX1042) );
and2 gate( .a(N3641), .b(p418), .O(EX1043) );
and2 gate( .a(N2646_NOT), .b(EX1043), .O(EX1044) );
and2 gate( .a(N3641_NOT), .b(p419), .O(EX1045) );
and2 gate( .a(N2646), .b(EX1045), .O(EX1046) );
and2 gate( .a(N3641), .b(p420), .O(EX1047) );
and2 gate( .a(N2646), .b(EX1047), .O(EX1048) );
or2  gate( .a(EX1042), .b(EX1044), .O(EX1049) );
or2  gate( .a(EX1046), .b(EX1049), .O(EX1050) );
or2  gate( .a(EX1048), .b(EX1050), .O(N3720) );
and2 gate1073( .a(N3644), .b(N3557), .O(N3721) );
or3 gate1074( .a(N3651), .b(N3652), .c(N3653), .O(N3731) );
and2 gate1075( .a(N3657), .b(N3568), .O(N3734) );
and2 gate1076( .a(N3661), .b(N3573), .O(N3740) );
and2 gate1077( .a(N3663), .b(N3578), .O(N3743) );
or3 gate1078( .a(N3670), .b(N3671), .c(N3672), .O(N3753) );
and2 gate1079( .a(N3676), .b(N3589), .O(N3756) );
and2 gate1080( .a(N3680), .b(N3594), .O(N3762) );
inv1 gate1081( .a(N3643), .O(N3765) );
inv1 gate1082( .a(N3662), .O(N3766) );
inv1 gate( .a(N3705),.O(N3705_NOT) );
inv1 gate( .a(N3706),.O(N3706_NOT));
and2 gate( .a(N3705_NOT), .b(p421), .O(EX1051) );
and2 gate( .a(N3706_NOT), .b(EX1051), .O(EX1052) );
and2 gate( .a(N3705), .b(p422), .O(EX1053) );
and2 gate( .a(N3706_NOT), .b(EX1053), .O(EX1054) );
and2 gate( .a(N3705_NOT), .b(p423), .O(EX1055) );
and2 gate( .a(N3706), .b(EX1055), .O(EX1056) );
and2 gate( .a(N3705), .b(p424), .O(EX1057) );
and2 gate( .a(N3706), .b(EX1057), .O(EX1058) );
or2  gate( .a(EX1052), .b(EX1054), .O(EX1059) );
or2  gate( .a(EX1056), .b(EX1059), .O(EX1060) );
or2  gate( .a(EX1058), .b(EX1060), .O(N3773) );
inv1 gate( .a(N3707),.O(N3707_NOT) );
inv1 gate( .a(N3708),.O(N3708_NOT));
and2 gate( .a(N3707_NOT), .b(p425), .O(EX1061) );
and2 gate( .a(N3708_NOT), .b(EX1061), .O(EX1062) );
and2 gate( .a(N3707), .b(p426), .O(EX1063) );
and2 gate( .a(N3708_NOT), .b(EX1063), .O(EX1064) );
and2 gate( .a(N3707_NOT), .b(p427), .O(EX1065) );
and2 gate( .a(N3708), .b(EX1065), .O(EX1066) );
and2 gate( .a(N3707), .b(p428), .O(EX1067) );
and2 gate( .a(N3708), .b(EX1067), .O(EX1068) );
or2  gate( .a(EX1062), .b(EX1064), .O(EX1069) );
or2  gate( .a(EX1066), .b(EX1069), .O(EX1070) );
or2  gate( .a(EX1068), .b(EX1070), .O(N3774) );
inv1 gate( .a(N3700),.O(N3700_NOT) );
inv1 gate( .a(N3628),.O(N3628_NOT));
and2 gate( .a(N3700_NOT), .b(p429), .O(EX1071) );
and2 gate( .a(N3628_NOT), .b(EX1071), .O(EX1072) );
and2 gate( .a(N3700), .b(p430), .O(EX1073) );
and2 gate( .a(N3628_NOT), .b(EX1073), .O(EX1074) );
and2 gate( .a(N3700_NOT), .b(p431), .O(EX1075) );
and2 gate( .a(N3628), .b(EX1075), .O(EX1076) );
and2 gate( .a(N3700), .b(p432), .O(EX1077) );
and2 gate( .a(N3628), .b(EX1077), .O(EX1078) );
or2  gate( .a(EX1072), .b(EX1074), .O(EX1079) );
or2  gate( .a(EX1076), .b(EX1079), .O(EX1080) );
or2  gate( .a(EX1078), .b(EX1080), .O(N3775) );
inv1 gate1086( .a(N3700), .O(N3776) );
nand2 gate1087( .a(N3697), .b(N3629), .O(N3777) );
inv1 gate1088( .a(N3697), .O(N3778) );
and2 gate1089( .a(N3712), .b(N2645), .O(N3779) );
and2 gate1090( .a(N3711), .b(N2647), .O(N3780) );
or2 gate1091( .a(N3645), .b(N3648), .O(N3786) );
nor2 gate1092( .a(N3645), .b(N3648), .O(N3789) );
or2 gate1093( .a(N3664), .b(N3667), .O(N3800) );
nor2 gate1094( .a(N3664), .b(N3667), .O(N3803) );
and2 gate1095( .a(N3654), .b(N1917), .O(N3809) );
and2 gate1096( .a(N3658), .b(N1917), .O(N3812) );
and2 gate1097( .a(N3673), .b(N1926), .O(N3815) );
inv1 gate( .a(N3677),.O(N3677_NOT) );
inv1 gate( .a(N1926),.O(N1926_NOT));
and2 gate( .a(N3677_NOT), .b(p433), .O(EX1081) );
and2 gate( .a(N1926_NOT), .b(EX1081), .O(EX1082) );
and2 gate( .a(N3677), .b(p434), .O(EX1083) );
and2 gate( .a(N1926_NOT), .b(EX1083), .O(EX1084) );
and2 gate( .a(N3677_NOT), .b(p435), .O(EX1085) );
and2 gate( .a(N1926), .b(EX1085), .O(EX1086) );
and2 gate( .a(N3677), .b(p436), .O(EX1087) );
and2 gate( .a(N1926), .b(EX1087), .O(EX1088) );
or2  gate( .a(EX1082), .b(EX1084), .O(EX1089) );
or2  gate( .a(EX1086), .b(EX1089), .O(EX1090) );
or2  gate( .a(EX1088), .b(EX1090), .O(N3818) );
buf1 gate1099( .a(N3682), .O(N3821) );
buf1 gate1100( .a(N3682), .O(N3824) );
buf1 gate1101( .a(N3690), .O(N3827) );
buf1 gate1102( .a(N3690), .O(N3830) );
nand2 gate1103( .a(N3773), .b(N3774), .O(N3833) );
inv1 gate( .a(N3487),.O(N3487_NOT) );
inv1 gate( .a(N3776),.O(N3776_NOT));
and2 gate( .a(N3487_NOT), .b(p437), .O(EX1091) );
and2 gate( .a(N3776_NOT), .b(EX1091), .O(EX1092) );
and2 gate( .a(N3487), .b(p438), .O(EX1093) );
and2 gate( .a(N3776_NOT), .b(EX1093), .O(EX1094) );
and2 gate( .a(N3487_NOT), .b(p439), .O(EX1095) );
and2 gate( .a(N3776), .b(EX1095), .O(EX1096) );
and2 gate( .a(N3487), .b(p440), .O(EX1097) );
and2 gate( .a(N3776), .b(EX1097), .O(EX1098) );
or2  gate( .a(EX1092), .b(EX1094), .O(EX1099) );
or2  gate( .a(EX1096), .b(EX1099), .O(EX1100) );
or2  gate( .a(EX1098), .b(EX1100), .O(N3834) );
nand2 gate1105( .a(N3484), .b(N3778), .O(N3835) );
and2 gate1106( .a(N3789), .b(N3731), .O(N3838) );
and2 gate1107( .a(N3803), .b(N3753), .O(N3845) );
buf1 gate1108( .a(N3721), .O(N3850) );
buf1 gate1109( .a(N3734), .O(N3855) );
buf1 gate1110( .a(N3740), .O(N3858) );
buf1 gate1111( .a(N3743), .O(N3861) );
buf1 gate1112( .a(N3756), .O(N3865) );
buf1 gate1113( .a(N3762), .O(N3868) );
nand2 gate1114( .a(N3775), .b(N3834), .O(N3884) );
nand2 gate1115( .a(N3777), .b(N3835), .O(N3885) );
nand2 gate1116( .a(N3721), .b(N3786), .O(N3894) );
nand2 gate1117( .a(N3743), .b(N3800), .O(N3895) );
inv1 gate1118( .a(N3821), .O(N3898) );
inv1 gate1119( .a(N3824), .O(N3899) );
inv1 gate1120( .a(N3830), .O(N3906) );
inv1 gate1121( .a(N3827), .O(N3911) );
and2 gate1122( .a(N3786), .b(N1912), .O(N3912) );
buf1 gate1123( .a(N3812), .O(N3913) );
and2 gate1124( .a(N3800), .b(N1917), .O(N3916) );
buf1 gate1125( .a(N3818), .O(N3917) );
inv1 gate1126( .a(N3809), .O(N3920) );
buf1 gate1127( .a(N3818), .O(N3921) );
inv1 gate1128( .a(N3884), .O(N3924) );
inv1 gate1129( .a(N3885), .O(N3925) );
and4 gate1130( .a(N3721), .b(N3838), .c(N3734), .d(N3740), .O(N3926) );
nand3 gate1131( .a(N3721), .b(N3838), .c(N3654), .O(N3930) );
nand4 gate1132( .a(N3658), .b(N3838), .c(N3734), .d(N3721), .O(N3931) );
and4 gate1133( .a(N3743), .b(N3845), .c(N3756), .d(N3762), .O(N3932) );
nand3 gate1134( .a(N3743), .b(N3845), .c(N3673), .O(N3935) );
nand4 gate1135( .a(N3677), .b(N3845), .c(N3756), .d(N3743), .O(N3936) );
buf1 gate1136( .a(N3838), .O(N3937) );
buf1 gate1137( .a(N3845), .O(N3940) );
inv1 gate1138( .a(N3912), .O(N3947) );
inv1 gate1139( .a(N3916), .O(N3948) );
buf1 gate1140( .a(N3850), .O(N3950) );
buf1 gate1141( .a(N3850), .O(N3953) );
buf1 gate1142( .a(N3855), .O(N3956) );
buf1 gate1143( .a(N3855), .O(N3959) );
buf1 gate1144( .a(N3858), .O(N3962) );
buf1 gate1145( .a(N3858), .O(N3965) );
buf1 gate1146( .a(N3861), .O(N3968) );
buf1 gate1147( .a(N3861), .O(N3971) );
buf1 gate1148( .a(N3865), .O(N3974) );
buf1 gate1149( .a(N3865), .O(N3977) );
buf1 gate1150( .a(N3868), .O(N3980) );
buf1 gate1151( .a(N3868), .O(N3983) );
nand2 gate1152( .a(N3924), .b(N3925), .O(N3987) );
nand4 gate1153( .a(N3765), .b(N3894), .c(N3930), .d(N3931), .O(N3992) );
nand4 gate1154( .a(N3766), .b(N3895), .c(N3935), .d(N3936), .O(N3996) );
inv1 gate1155( .a(N3921), .O(N4013) );
and2 gate1156( .a(N3932), .b(N3926), .O(N4028) );
nand2 gate1157( .a(N3953), .b(N3681), .O(N4029) );
nand2 gate1158( .a(N3959), .b(N3686), .O(N4030) );
nand2 gate1159( .a(N3965), .b(N3688), .O(N4031) );
nand2 gate1160( .a(N3971), .b(N3689), .O(N4032) );
nand2 gate1161( .a(N3977), .b(N3693), .O(N4033) );
nand2 gate1162( .a(N3983), .b(N3695), .O(N4034) );
buf1 gate1163( .a(N3926), .O(N4035) );
inv1 gate1164( .a(N3953), .O(N4042) );
inv1 gate1165( .a(N3956), .O(N4043) );
inv1 gate( .a(N3956),.O(N3956_NOT) );
inv1 gate( .a(N3685),.O(N3685_NOT));
and2 gate( .a(N3956_NOT), .b(p441), .O(EX1101) );
and2 gate( .a(N3685_NOT), .b(EX1101), .O(EX1102) );
and2 gate( .a(N3956), .b(p442), .O(EX1103) );
and2 gate( .a(N3685_NOT), .b(EX1103), .O(EX1104) );
and2 gate( .a(N3956_NOT), .b(p443), .O(EX1105) );
and2 gate( .a(N3685), .b(EX1105), .O(EX1106) );
and2 gate( .a(N3956), .b(p444), .O(EX1107) );
and2 gate( .a(N3685), .b(EX1107), .O(EX1108) );
or2  gate( .a(EX1102), .b(EX1104), .O(EX1109) );
or2  gate( .a(EX1106), .b(EX1109), .O(EX1110) );
or2  gate( .a(EX1108), .b(EX1110), .O(N4044) );
inv1 gate1167( .a(N3959), .O(N4045) );
inv1 gate1168( .a(N3962), .O(N4046) );
nand2 gate1169( .a(N3962), .b(N3687), .O(N4047) );
inv1 gate1170( .a(N3965), .O(N4048) );
inv1 gate1171( .a(N3971), .O(N4049) );
inv1 gate1172( .a(N3977), .O(N4050) );
inv1 gate1173( .a(N3980), .O(N4051) );
inv1 gate( .a(N3980),.O(N3980_NOT) );
inv1 gate( .a(N3694),.O(N3694_NOT));
and2 gate( .a(N3980_NOT), .b(p445), .O(EX1111) );
and2 gate( .a(N3694_NOT), .b(EX1111), .O(EX1112) );
and2 gate( .a(N3980), .b(p446), .O(EX1113) );
and2 gate( .a(N3694_NOT), .b(EX1113), .O(EX1114) );
and2 gate( .a(N3980_NOT), .b(p447), .O(EX1115) );
and2 gate( .a(N3694), .b(EX1115), .O(EX1116) );
and2 gate( .a(N3980), .b(p448), .O(EX1117) );
and2 gate( .a(N3694), .b(EX1117), .O(EX1118) );
or2  gate( .a(EX1112), .b(EX1114), .O(EX1119) );
or2  gate( .a(EX1116), .b(EX1119), .O(EX1120) );
or2  gate( .a(EX1118), .b(EX1120), .O(N4052) );
inv1 gate1175( .a(N3983), .O(N4053) );
inv1 gate1176( .a(N3974), .O(N4054) );
nand2 gate1177( .a(N3974), .b(N3696), .O(N4055) );
and2 gate1178( .a(N3932), .b(N2304), .O(N4056) );
inv1 gate1179( .a(N3950), .O(N4057) );
nand2 gate1180( .a(N3950), .b(N3703), .O(N4058) );
buf1 gate1181( .a(N3937), .O(N4059) );
buf1 gate1182( .a(N3937), .O(N4062) );
inv1 gate1183( .a(N3968), .O(N4065) );
nand2 gate1184( .a(N3968), .b(N3704), .O(N4066) );
buf1 gate1185( .a(N3940), .O(N4067) );
buf1 gate1186( .a(N3940), .O(N4070) );
nand2 gate1187( .a(N3926), .b(N3996), .O(N4073) );
inv1 gate1188( .a(N3992), .O(N4074) );
nand2 gate1189( .a(N3493), .b(N4042), .O(N4075) );
nand2 gate1190( .a(N3499), .b(N4045), .O(N4076) );
nand2 gate1191( .a(N3505), .b(N4048), .O(N4077) );
nand2 gate1192( .a(N3511), .b(N4049), .O(N4078) );
nand2 gate1193( .a(N3517), .b(N4050), .O(N4079) );
nand2 gate1194( .a(N3523), .b(N4053), .O(N4080) );
nand2 gate1195( .a(N3496), .b(N4043), .O(N4085) );
nand2 gate1196( .a(N3502), .b(N4046), .O(N4086) );
nand2 gate1197( .a(N3520), .b(N4051), .O(N4088) );
nand2 gate1198( .a(N3514), .b(N4054), .O(N4090) );
and2 gate1199( .a(N3996), .b(N1926), .O(N4091) );
or2 gate1200( .a(N3605), .b(N4056), .O(N4094) );
nand2 gate1201( .a(N3490), .b(N4057), .O(N4098) );
inv1 gate( .a(N3508),.O(N3508_NOT) );
inv1 gate( .a(N4065),.O(N4065_NOT));
and2 gate( .a(N3508_NOT), .b(p449), .O(EX1121) );
and2 gate( .a(N4065_NOT), .b(EX1121), .O(EX1122) );
and2 gate( .a(N3508), .b(p450), .O(EX1123) );
and2 gate( .a(N4065_NOT), .b(EX1123), .O(EX1124) );
and2 gate( .a(N3508_NOT), .b(p451), .O(EX1125) );
and2 gate( .a(N4065), .b(EX1125), .O(EX1126) );
and2 gate( .a(N3508), .b(p452), .O(EX1127) );
and2 gate( .a(N4065), .b(EX1127), .O(EX1128) );
or2  gate( .a(EX1122), .b(EX1124), .O(EX1129) );
or2  gate( .a(EX1126), .b(EX1129), .O(EX1130) );
or2  gate( .a(EX1128), .b(EX1130), .O(N4101) );
inv1 gate( .a(N4073),.O(N4073_NOT) );
inv1 gate( .a(N4074),.O(N4074_NOT));
and2 gate( .a(N4073_NOT), .b(p453), .O(EX1131) );
and2 gate( .a(N4074_NOT), .b(EX1131), .O(EX1132) );
and2 gate( .a(N4073), .b(p454), .O(EX1133) );
and2 gate( .a(N4074_NOT), .b(EX1133), .O(EX1134) );
and2 gate( .a(N4073_NOT), .b(p455), .O(EX1135) );
and2 gate( .a(N4074), .b(EX1135), .O(EX1136) );
and2 gate( .a(N4073), .b(p456), .O(EX1137) );
and2 gate( .a(N4074), .b(EX1137), .O(EX1138) );
or2  gate( .a(EX1132), .b(EX1134), .O(EX1139) );
or2  gate( .a(EX1136), .b(EX1139), .O(EX1140) );
or2  gate( .a(EX1138), .b(EX1140), .O(N4104) );
inv1 gate( .a(N4075),.O(N4075_NOT) );
inv1 gate( .a(N4029),.O(N4029_NOT));
and2 gate( .a(N4075_NOT), .b(p457), .O(EX1141) );
and2 gate( .a(N4029_NOT), .b(EX1141), .O(EX1142) );
and2 gate( .a(N4075), .b(p458), .O(EX1143) );
and2 gate( .a(N4029_NOT), .b(EX1143), .O(EX1144) );
and2 gate( .a(N4075_NOT), .b(p459), .O(EX1145) );
and2 gate( .a(N4029), .b(EX1145), .O(EX1146) );
and2 gate( .a(N4075), .b(p460), .O(EX1147) );
and2 gate( .a(N4029), .b(EX1147), .O(EX1148) );
or2  gate( .a(EX1142), .b(EX1144), .O(EX1149) );
or2  gate( .a(EX1146), .b(EX1149), .O(EX1150) );
or2  gate( .a(EX1148), .b(EX1150), .O(N4105) );
nand2 gate1205( .a(N4062), .b(N3899), .O(N4106) );
nand2 gate1206( .a(N4076), .b(N4030), .O(N4107) );
nand2 gate1207( .a(N4077), .b(N4031), .O(N4108) );
nand2 gate1208( .a(N4078), .b(N4032), .O(N4109) );
nand2 gate1209( .a(N4070), .b(N3906), .O(N4110) );
inv1 gate( .a(N4079),.O(N4079_NOT) );
inv1 gate( .a(N4033),.O(N4033_NOT));
and2 gate( .a(N4079_NOT), .b(p461), .O(EX1151) );
and2 gate( .a(N4033_NOT), .b(EX1151), .O(EX1152) );
and2 gate( .a(N4079), .b(p462), .O(EX1153) );
and2 gate( .a(N4033_NOT), .b(EX1153), .O(EX1154) );
and2 gate( .a(N4079_NOT), .b(p463), .O(EX1155) );
and2 gate( .a(N4033), .b(EX1155), .O(EX1156) );
and2 gate( .a(N4079), .b(p464), .O(EX1157) );
and2 gate( .a(N4033), .b(EX1157), .O(EX1158) );
or2  gate( .a(EX1152), .b(EX1154), .O(EX1159) );
or2  gate( .a(EX1156), .b(EX1159), .O(EX1160) );
or2  gate( .a(EX1158), .b(EX1160), .O(N4111) );
nand2 gate1211( .a(N4080), .b(N4034), .O(N4112) );
inv1 gate1212( .a(N4059), .O(N4113) );
nand2 gate1213( .a(N4059), .b(N3898), .O(N4114) );
inv1 gate1214( .a(N4062), .O(N4115) );
nand2 gate1215( .a(N4085), .b(N4044), .O(N4116) );
nand2 gate1216( .a(N4086), .b(N4047), .O(N4119) );
inv1 gate1217( .a(N4070), .O(N4122) );
nand2 gate1218( .a(N4088), .b(N4052), .O(N4123) );
inv1 gate1219( .a(N4067), .O(N4126) );
nand2 gate1220( .a(N4067), .b(N3911), .O(N4127) );
inv1 gate( .a(N4090),.O(N4090_NOT) );
inv1 gate( .a(N4055),.O(N4055_NOT));
and2 gate( .a(N4090_NOT), .b(p465), .O(EX1161) );
and2 gate( .a(N4055_NOT), .b(EX1161), .O(EX1162) );
and2 gate( .a(N4090), .b(p466), .O(EX1163) );
and2 gate( .a(N4055_NOT), .b(EX1163), .O(EX1164) );
and2 gate( .a(N4090_NOT), .b(p467), .O(EX1165) );
and2 gate( .a(N4055), .b(EX1165), .O(EX1166) );
and2 gate( .a(N4090), .b(p468), .O(EX1167) );
and2 gate( .a(N4055), .b(EX1167), .O(EX1168) );
or2  gate( .a(EX1162), .b(EX1164), .O(EX1169) );
or2  gate( .a(EX1166), .b(EX1169), .O(EX1170) );
or2  gate( .a(EX1168), .b(EX1170), .O(N4128) );
nand2 gate1222( .a(N4098), .b(N4058), .O(N4139) );
nand2 gate1223( .a(N4101), .b(N4066), .O(N4142) );
inv1 gate1224( .a(N4104), .O(N4145) );
inv1 gate1225( .a(N4105), .O(N4146) );
inv1 gate( .a(N3824),.O(N3824_NOT) );
inv1 gate( .a(N4115),.O(N4115_NOT));
and2 gate( .a(N3824_NOT), .b(p469), .O(EX1171) );
and2 gate( .a(N4115_NOT), .b(EX1171), .O(EX1172) );
and2 gate( .a(N3824), .b(p470), .O(EX1173) );
and2 gate( .a(N4115_NOT), .b(EX1173), .O(EX1174) );
and2 gate( .a(N3824_NOT), .b(p471), .O(EX1175) );
and2 gate( .a(N4115), .b(EX1175), .O(EX1176) );
and2 gate( .a(N3824), .b(p472), .O(EX1177) );
and2 gate( .a(N4115), .b(EX1177), .O(EX1178) );
or2  gate( .a(EX1172), .b(EX1174), .O(EX1179) );
or2  gate( .a(EX1176), .b(EX1179), .O(EX1180) );
or2  gate( .a(EX1178), .b(EX1180), .O(N4147) );
inv1 gate1227( .a(N4107), .O(N4148) );
inv1 gate1228( .a(N4108), .O(N4149) );
inv1 gate1229( .a(N4109), .O(N4150) );
nand2 gate1230( .a(N3830), .b(N4122), .O(N4151) );
inv1 gate1231( .a(N4111), .O(N4152) );
inv1 gate1232( .a(N4112), .O(N4153) );
nand2 gate1233( .a(N3821), .b(N4113), .O(N4154) );
nand2 gate1234( .a(N3827), .b(N4126), .O(N4161) );
buf1 gate1235( .a(N4091), .O(N4167) );
buf1 gate1236( .a(N4094), .O(N4174) );
buf1 gate1237( .a(N4091), .O(N4182) );
and2 gate1238( .a(N330), .b(N4094), .O(N4186) );
and2 gate1239( .a(N4146), .b(N2230), .O(N4189) );
nand2 gate1240( .a(N4147), .b(N4106), .O(N4190) );
inv1 gate( .a(N4148),.O(N4148_NOT) );
inv1 gate( .a(N2232),.O(N2232_NOT));
and2 gate( .a(N4148_NOT), .b(p473), .O(EX1181) );
and2 gate( .a(N2232_NOT), .b(EX1181), .O(EX1182) );
and2 gate( .a(N4148), .b(p474), .O(EX1183) );
and2 gate( .a(N2232_NOT), .b(EX1183), .O(EX1184) );
and2 gate( .a(N4148_NOT), .b(p475), .O(EX1185) );
and2 gate( .a(N2232), .b(EX1185), .O(EX1186) );
and2 gate( .a(N4148), .b(p476), .O(EX1187) );
and2 gate( .a(N2232), .b(EX1187), .O(EX1188) );
or2  gate( .a(EX1182), .b(EX1184), .O(EX1189) );
or2  gate( .a(EX1186), .b(EX1189), .O(EX1190) );
or2  gate( .a(EX1188), .b(EX1190), .O(N4191) );
and2 gate1242( .a(N4149), .b(N2233), .O(N4192) );
and2 gate1243( .a(N4150), .b(N2234), .O(N4193) );
nand2 gate1244( .a(N4151), .b(N4110), .O(N4194) );
and2 gate1245( .a(N4152), .b(N2236), .O(N4195) );
and2 gate1246( .a(N4153), .b(N2237), .O(N4196) );
nand2 gate1247( .a(N4154), .b(N4114), .O(N4197) );
buf1 gate1248( .a(N4116), .O(N4200) );
buf1 gate1249( .a(N4116), .O(N4203) );
buf1 gate1250( .a(N4119), .O(N4209) );
buf1 gate1251( .a(N4119), .O(N4213) );
inv1 gate( .a(N4161),.O(N4161_NOT) );
inv1 gate( .a(N4127),.O(N4127_NOT));
and2 gate( .a(N4161_NOT), .b(p477), .O(EX1191) );
and2 gate( .a(N4127_NOT), .b(EX1191), .O(EX1192) );
and2 gate( .a(N4161), .b(p478), .O(EX1193) );
and2 gate( .a(N4127_NOT), .b(EX1193), .O(EX1194) );
and2 gate( .a(N4161_NOT), .b(p479), .O(EX1195) );
and2 gate( .a(N4127), .b(EX1195), .O(EX1196) );
and2 gate( .a(N4161), .b(p480), .O(EX1197) );
and2 gate( .a(N4127), .b(EX1197), .O(EX1198) );
or2  gate( .a(EX1192), .b(EX1194), .O(EX1199) );
or2  gate( .a(EX1196), .b(EX1199), .O(EX1200) );
or2  gate( .a(EX1198), .b(EX1200), .O(N4218) );
buf1 gate1253( .a(N4123), .O(N4223) );
and2 gate1254( .a(N4128), .b(N3917), .O(N4238) );
inv1 gate1255( .a(N4139), .O(N4239) );
inv1 gate1256( .a(N4142), .O(N4241) );
and2 gate1257( .a(N330), .b(N4123), .O(N4242) );
buf1 gate1258( .a(N4128), .O(N4247) );
nor3 gate1259( .a(N3713), .b(N4189), .c(N2898), .O(N4251) );
inv1 gate1260( .a(N4190), .O(N4252) );
nor3 gate1261( .a(N3715), .b(N4191), .c(N2900), .O(N4253) );
nor3 gate1262( .a(N3716), .b(N4192), .c(N2901), .O(N4254) );
nor3 gate1263( .a(N3717), .b(N4193), .c(N3406), .O(N4255) );
inv1 gate1264( .a(N4194), .O(N4256) );
nor3 gate1265( .a(N3719), .b(N4195), .c(N3779), .O(N4257) );
nor3 gate1266( .a(N3720), .b(N4196), .c(N3780), .O(N4258) );
and2 gate1267( .a(N4167), .b(N4035), .O(N4283) );
inv1 gate( .a(N4174),.O(N4174_NOT) );
inv1 gate( .a(N4035),.O(N4035_NOT));
and2 gate( .a(N4174_NOT), .b(p481), .O(EX1201) );
and2 gate( .a(N4035_NOT), .b(EX1201), .O(EX1202) );
and2 gate( .a(N4174), .b(p482), .O(EX1203) );
and2 gate( .a(N4035_NOT), .b(EX1203), .O(EX1204) );
and2 gate( .a(N4174_NOT), .b(p483), .O(EX1205) );
and2 gate( .a(N4035), .b(EX1205), .O(EX1206) );
and2 gate( .a(N4174), .b(p484), .O(EX1207) );
and2 gate( .a(N4035), .b(EX1207), .O(EX1208) );
or2  gate( .a(EX1202), .b(EX1204), .O(EX1209) );
or2  gate( .a(EX1206), .b(EX1209), .O(EX1210) );
or2  gate( .a(EX1208), .b(EX1210), .O(N4284) );
or2 gate1269( .a(N3815), .b(N4238), .O(N4287) );
inv1 gate1270( .a(N4186), .O(N4291) );
inv1 gate1271( .a(N4167), .O(N4295) );
buf1 gate1272( .a(N4167), .O(N4296) );
inv1 gate1273( .a(N4182), .O(N4299) );
and2 gate1274( .a(N4252), .b(N2231), .O(N4303) );
and2 gate1275( .a(N4256), .b(N2235), .O(N4304) );
buf1 gate1276( .a(N4197), .O(N4305) );
inv1 gate( .a(N3992),.O(N3992_NOT) );
inv1 gate( .a(N4283),.O(N4283_NOT));
and2 gate( .a(N3992_NOT), .b(p485), .O(EX1211) );
and2 gate( .a(N4283_NOT), .b(EX1211), .O(EX1212) );
and2 gate( .a(N3992), .b(p486), .O(EX1213) );
and2 gate( .a(N4283_NOT), .b(EX1213), .O(EX1214) );
and2 gate( .a(N3992_NOT), .b(p487), .O(EX1215) );
and2 gate( .a(N4283), .b(EX1215), .O(EX1216) );
and2 gate( .a(N3992), .b(p488), .O(EX1217) );
and2 gate( .a(N4283), .b(EX1217), .O(EX1218) );
or2  gate( .a(EX1212), .b(EX1214), .O(EX1219) );
or2  gate( .a(EX1216), .b(EX1219), .O(EX1220) );
or2  gate( .a(EX1218), .b(EX1220), .O(N4310) );
and3 gate1278( .a(N4174), .b(N4213), .c(N4203), .O(N4316) );
and2 gate1279( .a(N4174), .b(N4209), .O(N4317) );
and3 gate1280( .a(N4223), .b(N4128), .c(N4218), .O(N4318) );
and2 gate1281( .a(N4223), .b(N4128), .O(N4319) );
and2 gate1282( .a(N4167), .b(N4209), .O(N4322) );
nand2 gate1283( .a(N4203), .b(N3913), .O(N4325) );
nand3 gate1284( .a(N4203), .b(N4213), .c(N4167), .O(N4326) );
nand2 gate1285( .a(N4218), .b(N3815), .O(N4327) );
nand3 gate1286( .a(N4218), .b(N4128), .c(N3917), .O(N4328) );
nand2 gate1287( .a(N4247), .b(N4013), .O(N4329) );
inv1 gate1288( .a(N4247), .O(N4330) );
and3 gate1289( .a(N330), .b(N4094), .c(N4295), .O(N4331) );
inv1 gate( .a(N4251),.O(N4251_NOT) );
inv1 gate( .a(N2730),.O(N2730_NOT));
and2 gate( .a(N4251_NOT), .b(p489), .O(EX1221) );
and2 gate( .a(N2730_NOT), .b(EX1221), .O(EX1222) );
and2 gate( .a(N4251), .b(p490), .O(EX1223) );
and2 gate( .a(N2730_NOT), .b(EX1223), .O(EX1224) );
and2 gate( .a(N4251_NOT), .b(p491), .O(EX1225) );
and2 gate( .a(N2730), .b(EX1225), .O(EX1226) );
and2 gate( .a(N4251), .b(p492), .O(EX1227) );
and2 gate( .a(N2730), .b(EX1227), .O(EX1228) );
or2  gate( .a(EX1222), .b(EX1224), .O(EX1229) );
or2  gate( .a(EX1226), .b(EX1229), .O(EX1230) );
or2  gate( .a(EX1228), .b(EX1230), .O(N4335) );
inv1 gate( .a(N4253),.O(N4253_NOT) );
inv1 gate( .a(N2734),.O(N2734_NOT));
and2 gate( .a(N4253_NOT), .b(p493), .O(EX1231) );
and2 gate( .a(N2734_NOT), .b(EX1231), .O(EX1232) );
and2 gate( .a(N4253), .b(p494), .O(EX1233) );
and2 gate( .a(N2734_NOT), .b(EX1233), .O(EX1234) );
and2 gate( .a(N4253_NOT), .b(p495), .O(EX1235) );
and2 gate( .a(N2734), .b(EX1235), .O(EX1236) );
and2 gate( .a(N4253), .b(p496), .O(EX1237) );
and2 gate( .a(N2734), .b(EX1237), .O(EX1238) );
or2  gate( .a(EX1232), .b(EX1234), .O(EX1239) );
or2  gate( .a(EX1236), .b(EX1239), .O(EX1240) );
or2  gate( .a(EX1238), .b(EX1240), .O(N4338) );
inv1 gate( .a(N4254),.O(N4254_NOT) );
inv1 gate( .a(N2736),.O(N2736_NOT));
and2 gate( .a(N4254_NOT), .b(p497), .O(EX1241) );
and2 gate( .a(N2736_NOT), .b(EX1241), .O(EX1242) );
and2 gate( .a(N4254), .b(p498), .O(EX1243) );
and2 gate( .a(N2736_NOT), .b(EX1243), .O(EX1244) );
and2 gate( .a(N4254_NOT), .b(p499), .O(EX1245) );
and2 gate( .a(N2736), .b(EX1245), .O(EX1246) );
and2 gate( .a(N4254), .b(p500), .O(EX1247) );
and2 gate( .a(N2736), .b(EX1247), .O(EX1248) );
or2  gate( .a(EX1242), .b(EX1244), .O(EX1249) );
or2  gate( .a(EX1246), .b(EX1249), .O(EX1250) );
or2  gate( .a(EX1248), .b(EX1250), .O(N4341) );
inv1 gate( .a(N4255),.O(N4255_NOT) );
inv1 gate( .a(N2738),.O(N2738_NOT));
and2 gate( .a(N4255_NOT), .b(p501), .O(EX1251) );
and2 gate( .a(N2738_NOT), .b(EX1251), .O(EX1252) );
and2 gate( .a(N4255), .b(p502), .O(EX1253) );
and2 gate( .a(N2738_NOT), .b(EX1253), .O(EX1254) );
and2 gate( .a(N4255_NOT), .b(p503), .O(EX1255) );
and2 gate( .a(N2738), .b(EX1255), .O(EX1256) );
and2 gate( .a(N4255), .b(p504), .O(EX1257) );
and2 gate( .a(N2738), .b(EX1257), .O(EX1258) );
or2  gate( .a(EX1252), .b(EX1254), .O(EX1259) );
or2  gate( .a(EX1256), .b(EX1259), .O(EX1260) );
or2  gate( .a(EX1258), .b(EX1260), .O(N4344) );
and2 gate1294( .a(N4257), .b(N2742), .O(N4347) );
inv1 gate( .a(N4258),.O(N4258_NOT) );
inv1 gate( .a(N2744),.O(N2744_NOT));
and2 gate( .a(N4258_NOT), .b(p505), .O(EX1261) );
and2 gate( .a(N2744_NOT), .b(EX1261), .O(EX1262) );
and2 gate( .a(N4258), .b(p506), .O(EX1263) );
and2 gate( .a(N2744_NOT), .b(EX1263), .O(EX1264) );
and2 gate( .a(N4258_NOT), .b(p507), .O(EX1265) );
and2 gate( .a(N2744), .b(EX1265), .O(EX1266) );
and2 gate( .a(N4258), .b(p508), .O(EX1267) );
and2 gate( .a(N2744), .b(EX1267), .O(EX1268) );
or2  gate( .a(EX1262), .b(EX1264), .O(EX1269) );
or2  gate( .a(EX1266), .b(EX1269), .O(EX1270) );
or2  gate( .a(EX1268), .b(EX1270), .O(N4350) );
buf1 gate1296( .a(N4197), .O(N4353) );
buf1 gate1297( .a(N4203), .O(N4356) );
buf1 gate1298( .a(N4209), .O(N4359) );
buf1 gate1299( .a(N4218), .O(N4362) );
buf1 gate1300( .a(N4242), .O(N4365) );
buf1 gate1301( .a(N4242), .O(N4368) );
and2 gate1302( .a(N4223), .b(N4223), .O(N4371) );
nor3 gate1303( .a(N3714), .b(N4303), .c(N2899), .O(N4376) );
nor3 gate1304( .a(N3718), .b(N4304), .c(N3642), .O(N4377) );
and2 gate1305( .a(N330), .b(N4317), .O(N4387) );
and2 gate1306( .a(N330), .b(N4318), .O(N4390) );
nand2 gate1307( .a(N3921), .b(N4330), .O(N4393) );
buf1 gate1308( .a(N4287), .O(N4398) );
buf1 gate1309( .a(N4284), .O(N4413) );
nand3 gate1310( .a(N3920), .b(N4325), .c(N4326), .O(N4416) );
or2 gate1311( .a(N3812), .b(N4322), .O(N4421) );
nand3 gate1312( .a(N3948), .b(N4327), .c(N4328), .O(N4427) );
buf1 gate1313( .a(N4287), .O(N4430) );
inv1 gate( .a(N330),.O(N330_NOT) );
inv1 gate( .a(N4316),.O(N4316_NOT));
and2 gate( .a(N330_NOT), .b(p509), .O(EX1271) );
and2 gate( .a(N4316_NOT), .b(EX1271), .O(EX1272) );
and2 gate( .a(N330), .b(p510), .O(EX1273) );
and2 gate( .a(N4316_NOT), .b(EX1273), .O(EX1274) );
and2 gate( .a(N330_NOT), .b(p511), .O(EX1275) );
and2 gate( .a(N4316), .b(EX1275), .O(EX1276) );
and2 gate( .a(N330), .b(p512), .O(EX1277) );
and2 gate( .a(N4316), .b(EX1277), .O(EX1278) );
or2  gate( .a(EX1272), .b(EX1274), .O(EX1279) );
or2  gate( .a(EX1276), .b(EX1279), .O(EX1280) );
or2  gate( .a(EX1278), .b(EX1280), .O(N4435) );
or2 gate1315( .a(N4331), .b(N4296), .O(N4442) );
and4 gate1316( .a(N4174), .b(N4305), .c(N4203), .d(N4213), .O(N4443) );
nand2 gate1317( .a(N4305), .b(N3809), .O(N4446) );
nand3 gate1318( .a(N4305), .b(N4200), .c(N3913), .O(N4447) );
nand4 gate1319( .a(N4305), .b(N4200), .c(N4213), .d(N4167), .O(N4448) );
inv1 gate1320( .a(N4356), .O(N4452) );
nand2 gate1321( .a(N4329), .b(N4393), .O(N4458) );
inv1 gate1322( .a(N4365), .O(N4461) );
inv1 gate1323( .a(N4368), .O(N4462) );
nand2 gate1324( .a(N4371), .b(N1460), .O(N4463) );
inv1 gate1325( .a(N4371), .O(N4464) );
buf1 gate1326( .a(N4310), .O(N4465) );
nor2 gate1327( .a(N4331), .b(N4296), .O(N4468) );
and2 gate1328( .a(N4376), .b(N2732), .O(N4472) );
inv1 gate( .a(N4377),.O(N4377_NOT) );
inv1 gate( .a(N2740),.O(N2740_NOT));
and2 gate( .a(N4377_NOT), .b(p513), .O(EX1281) );
and2 gate( .a(N2740_NOT), .b(EX1281), .O(EX1282) );
and2 gate( .a(N4377), .b(p514), .O(EX1283) );
and2 gate( .a(N2740_NOT), .b(EX1283), .O(EX1284) );
and2 gate( .a(N4377_NOT), .b(p515), .O(EX1285) );
and2 gate( .a(N2740), .b(EX1285), .O(EX1286) );
and2 gate( .a(N4377), .b(p516), .O(EX1287) );
and2 gate( .a(N2740), .b(EX1287), .O(EX1288) );
or2  gate( .a(EX1282), .b(EX1284), .O(EX1289) );
or2  gate( .a(EX1286), .b(EX1289), .O(EX1290) );
or2  gate( .a(EX1288), .b(EX1290), .O(N4475) );
buf1 gate1330( .a(N4310), .O(N4479) );
inv1 gate1331( .a(N4353), .O(N4484) );
inv1 gate1332( .a(N4359), .O(N4486) );
nand2 gate1333( .a(N4359), .b(N4299), .O(N4487) );
inv1 gate1334( .a(N4362), .O(N4491) );
and2 gate1335( .a(N330), .b(N4319), .O(N4493) );
inv1 gate1336( .a(N4398), .O(N4496) );
and2 gate1337( .a(N4287), .b(N4398), .O(N4497) );
and2 gate1338( .a(N4442), .b(N1769), .O(N4498) );
nand4 gate1339( .a(N3947), .b(N4446), .c(N4447), .d(N4448), .O(N4503) );
inv1 gate1340( .a(N4413), .O(N4506) );
inv1 gate1341( .a(N4435), .O(N4507) );
inv1 gate1342( .a(N4421), .O(N4508) );
nand2 gate1343( .a(N4421), .b(N4452), .O(N4509) );
inv1 gate1344( .a(N4427), .O(N4510) );
inv1 gate( .a(N4427),.O(N4427_NOT) );
inv1 gate( .a(N4241),.O(N4241_NOT));
and2 gate( .a(N4427_NOT), .b(p517), .O(EX1291) );
and2 gate( .a(N4241_NOT), .b(EX1291), .O(EX1292) );
and2 gate( .a(N4427), .b(p518), .O(EX1293) );
and2 gate( .a(N4241_NOT), .b(EX1293), .O(EX1294) );
and2 gate( .a(N4427_NOT), .b(p519), .O(EX1295) );
and2 gate( .a(N4241), .b(EX1295), .O(EX1296) );
and2 gate( .a(N4427), .b(p520), .O(EX1297) );
and2 gate( .a(N4241), .b(EX1297), .O(EX1298) );
or2  gate( .a(EX1292), .b(EX1294), .O(EX1299) );
or2  gate( .a(EX1296), .b(EX1299), .O(EX1300) );
or2  gate( .a(EX1298), .b(EX1300), .O(N4511) );
inv1 gate( .a(N965),.O(N965_NOT) );
inv1 gate( .a(N4464),.O(N4464_NOT));
and2 gate( .a(N965_NOT), .b(p521), .O(EX1301) );
and2 gate( .a(N4464_NOT), .b(EX1301), .O(EX1302) );
and2 gate( .a(N965), .b(p522), .O(EX1303) );
and2 gate( .a(N4464_NOT), .b(EX1303), .O(EX1304) );
and2 gate( .a(N965_NOT), .b(p523), .O(EX1305) );
and2 gate( .a(N4464), .b(EX1305), .O(EX1306) );
and2 gate( .a(N965), .b(p524), .O(EX1307) );
and2 gate( .a(N4464), .b(EX1307), .O(EX1308) );
or2  gate( .a(EX1302), .b(EX1304), .O(EX1309) );
or2  gate( .a(EX1306), .b(EX1309), .O(EX1310) );
or2  gate( .a(EX1308), .b(EX1310), .O(N4515) );
inv1 gate1347( .a(N4416), .O(N4526) );
nand2 gate1348( .a(N4416), .b(N4484), .O(N4527) );
nand2 gate1349( .a(N4182), .b(N4486), .O(N4528) );
inv1 gate1350( .a(N4430), .O(N4529) );
nand2 gate1351( .a(N4430), .b(N4491), .O(N4530) );
buf1 gate1352( .a(N4387), .O(N4531) );
buf1 gate1353( .a(N4387), .O(N4534) );
buf1 gate1354( .a(N4390), .O(N4537) );
buf1 gate1355( .a(N4390), .O(N4540) );
and3 gate1356( .a(N330), .b(N4319), .c(N4496), .O(N4545) );
inv1 gate( .a(N330),.O(N330_NOT) );
inv1 gate( .a(N4443),.O(N4443_NOT));
and2 gate( .a(N330_NOT), .b(p525), .O(EX1311) );
and2 gate( .a(N4443_NOT), .b(EX1311), .O(EX1312) );
and2 gate( .a(N330), .b(p526), .O(EX1313) );
and2 gate( .a(N4443_NOT), .b(EX1313), .O(EX1314) );
and2 gate( .a(N330_NOT), .b(p527), .O(EX1315) );
and2 gate( .a(N4443), .b(EX1315), .O(EX1316) );
and2 gate( .a(N330), .b(p528), .O(EX1317) );
and2 gate( .a(N4443), .b(EX1317), .O(EX1318) );
or2  gate( .a(EX1312), .b(EX1314), .O(EX1319) );
or2  gate( .a(EX1316), .b(EX1319), .O(EX1320) );
or2  gate( .a(EX1318), .b(EX1320), .O(N4549) );
nand2 gate1358( .a(N4356), .b(N4508), .O(N4552) );
nand2 gate1359( .a(N4142), .b(N4510), .O(N4555) );
inv1 gate1360( .a(N4493), .O(N4558) );
nand2 gate1361( .a(N4463), .b(N4515), .O(N4559) );
inv1 gate1362( .a(N4465), .O(N4562) );
inv1 gate( .a(N4310),.O(N4310_NOT) );
inv1 gate( .a(N4465),.O(N4465_NOT));
and2 gate( .a(N4310_NOT), .b(p529), .O(EX1321) );
and2 gate( .a(N4465_NOT), .b(EX1321), .O(EX1322) );
and2 gate( .a(N4310), .b(p530), .O(EX1323) );
and2 gate( .a(N4465_NOT), .b(EX1323), .O(EX1324) );
and2 gate( .a(N4310_NOT), .b(p531), .O(EX1325) );
and2 gate( .a(N4465), .b(EX1325), .O(EX1326) );
and2 gate( .a(N4310), .b(p532), .O(EX1327) );
and2 gate( .a(N4465), .b(EX1327), .O(EX1328) );
or2  gate( .a(EX1322), .b(EX1324), .O(EX1329) );
or2  gate( .a(EX1326), .b(EX1329), .O(EX1330) );
or2  gate( .a(EX1328), .b(EX1330), .O(N4563) );
buf1 gate1364( .a(N4468), .O(N4564) );
inv1 gate1365( .a(N4479), .O(N4568) );
buf1 gate1366( .a(N4443), .O(N4569) );
nand2 gate1367( .a(N4353), .b(N4526), .O(N4572) );
inv1 gate( .a(N4362),.O(N4362_NOT) );
inv1 gate( .a(N4529),.O(N4529_NOT));
and2 gate( .a(N4362_NOT), .b(p533), .O(EX1331) );
and2 gate( .a(N4529_NOT), .b(EX1331), .O(EX1332) );
and2 gate( .a(N4362), .b(p534), .O(EX1333) );
and2 gate( .a(N4529_NOT), .b(EX1333), .O(EX1334) );
and2 gate( .a(N4362_NOT), .b(p535), .O(EX1335) );
and2 gate( .a(N4529), .b(EX1335), .O(EX1336) );
and2 gate( .a(N4362), .b(p536), .O(EX1337) );
and2 gate( .a(N4529), .b(EX1337), .O(EX1338) );
or2  gate( .a(EX1332), .b(EX1334), .O(EX1339) );
or2  gate( .a(EX1336), .b(EX1339), .O(EX1340) );
or2  gate( .a(EX1338), .b(EX1340), .O(N4573) );
nand2 gate1369( .a(N4487), .b(N4528), .O(N4576) );
buf1 gate1370( .a(N4458), .O(N4581) );
buf1 gate1371( .a(N4458), .O(N4584) );
or3 gate1372( .a(N2758), .b(N4498), .c(N2761), .O(N4587) );
nor3 gate1373( .a(N2758), .b(N4498), .c(N2761), .O(N4588) );
or2 gate1374( .a(N4545), .b(N4497), .O(N4589) );
nand2 gate1375( .a(N4552), .b(N4509), .O(N4593) );
inv1 gate1376( .a(N4531), .O(N4596) );
inv1 gate1377( .a(N4534), .O(N4597) );
nand2 gate1378( .a(N4555), .b(N4511), .O(N4599) );
inv1 gate1379( .a(N4537), .O(N4602) );
inv1 gate1380( .a(N4540), .O(N4603) );
and3 gate1381( .a(N330), .b(N4284), .c(N4562), .O(N4608) );
buf1 gate1382( .a(N4503), .O(N4613) );
buf1 gate1383( .a(N4503), .O(N4616) );
nand2 gate1384( .a(N4572), .b(N4527), .O(N4619) );
nand2 gate1385( .a(N4573), .b(N4530), .O(N4623) );
inv1 gate1386( .a(N4588), .O(N4628) );
nand2 gate1387( .a(N4569), .b(N4506), .O(N4629) );
inv1 gate1388( .a(N4569), .O(N4630) );
inv1 gate1389( .a(N4576), .O(N4635) );
nand2 gate1390( .a(N4576), .b(N4291), .O(N4636) );
inv1 gate1391( .a(N4581), .O(N4640) );
nand2 gate1392( .a(N4581), .b(N4461), .O(N4641) );
inv1 gate1393( .a(N4584), .O(N4642) );
nand2 gate1394( .a(N4584), .b(N4462), .O(N4643) );
nor2 gate1395( .a(N4608), .b(N4563), .O(N4644) );
inv1 gate( .a(N4559),.O(N4559_NOT) );
inv1 gate( .a(N2128),.O(N2128_NOT));
and2 gate( .a(N4559_NOT), .b(p537), .O(EX1341) );
and2 gate( .a(N2128_NOT), .b(EX1341), .O(EX1342) );
and2 gate( .a(N4559), .b(p538), .O(EX1343) );
and2 gate( .a(N2128_NOT), .b(EX1343), .O(EX1344) );
and2 gate( .a(N4559_NOT), .b(p539), .O(EX1345) );
and2 gate( .a(N2128), .b(EX1345), .O(EX1346) );
and2 gate( .a(N4559), .b(p540), .O(EX1347) );
and2 gate( .a(N2128), .b(EX1347), .O(EX1348) );
or2  gate( .a(EX1342), .b(EX1344), .O(EX1349) );
or2  gate( .a(EX1346), .b(EX1349), .O(EX1350) );
or2  gate( .a(EX1348), .b(EX1350), .O(N4647) );
and2 gate1397( .a(N4559), .b(N2743), .O(N4650) );
buf1 gate1398( .a(N4549), .O(N4656) );
buf1 gate1399( .a(N4549), .O(N4659) );
buf1 gate1400( .a(N4564), .O(N4664) );
and2 gate1401( .a(N4587), .b(N4628), .O(N4667) );
nand2 gate1402( .a(N4413), .b(N4630), .O(N4668) );
inv1 gate1403( .a(N4616), .O(N4669) );
inv1 gate( .a(N4616),.O(N4616_NOT) );
inv1 gate( .a(N4239),.O(N4239_NOT));
and2 gate( .a(N4616_NOT), .b(p541), .O(EX1351) );
and2 gate( .a(N4239_NOT), .b(EX1351), .O(EX1352) );
and2 gate( .a(N4616), .b(p542), .O(EX1353) );
and2 gate( .a(N4239_NOT), .b(EX1353), .O(EX1354) );
and2 gate( .a(N4616_NOT), .b(p543), .O(EX1355) );
and2 gate( .a(N4239), .b(EX1355), .O(EX1356) );
and2 gate( .a(N4616), .b(p544), .O(EX1357) );
and2 gate( .a(N4239), .b(EX1357), .O(EX1358) );
or2  gate( .a(EX1352), .b(EX1354), .O(EX1359) );
or2  gate( .a(EX1356), .b(EX1359), .O(EX1360) );
or2  gate( .a(EX1358), .b(EX1360), .O(N4670) );
inv1 gate1405( .a(N4619), .O(N4673) );
nand2 gate1406( .a(N4619), .b(N4507), .O(N4674) );
inv1 gate( .a(N4186),.O(N4186_NOT) );
inv1 gate( .a(N4635),.O(N4635_NOT));
and2 gate( .a(N4186_NOT), .b(p545), .O(EX1361) );
and2 gate( .a(N4635_NOT), .b(EX1361), .O(EX1362) );
and2 gate( .a(N4186), .b(p546), .O(EX1363) );
and2 gate( .a(N4635_NOT), .b(EX1363), .O(EX1364) );
and2 gate( .a(N4186_NOT), .b(p547), .O(EX1365) );
and2 gate( .a(N4635), .b(EX1365), .O(EX1366) );
and2 gate( .a(N4186), .b(p548), .O(EX1367) );
and2 gate( .a(N4635), .b(EX1367), .O(EX1368) );
or2  gate( .a(EX1362), .b(EX1364), .O(EX1369) );
or2  gate( .a(EX1366), .b(EX1369), .O(EX1370) );
or2  gate( .a(EX1368), .b(EX1370), .O(N4675) );
inv1 gate1408( .a(N4623), .O(N4676) );
nand2 gate1409( .a(N4623), .b(N4558), .O(N4677) );
inv1 gate( .a(N4365),.O(N4365_NOT) );
inv1 gate( .a(N4640),.O(N4640_NOT));
and2 gate( .a(N4365_NOT), .b(p549), .O(EX1371) );
and2 gate( .a(N4640_NOT), .b(EX1371), .O(EX1372) );
and2 gate( .a(N4365), .b(p550), .O(EX1373) );
and2 gate( .a(N4640_NOT), .b(EX1373), .O(EX1374) );
and2 gate( .a(N4365_NOT), .b(p551), .O(EX1375) );
and2 gate( .a(N4640), .b(EX1375), .O(EX1376) );
and2 gate( .a(N4365), .b(p552), .O(EX1377) );
and2 gate( .a(N4640), .b(EX1377), .O(EX1378) );
or2  gate( .a(EX1372), .b(EX1374), .O(EX1379) );
or2  gate( .a(EX1376), .b(EX1379), .O(EX1380) );
or2  gate( .a(EX1378), .b(EX1380), .O(N4678) );
nand2 gate1411( .a(N4368), .b(N4642), .O(N4679) );
inv1 gate1412( .a(N4613), .O(N4687) );
nand2 gate1413( .a(N4613), .b(N4568), .O(N4688) );
buf1 gate1414( .a(N4593), .O(N4691) );
buf1 gate1415( .a(N4593), .O(N4694) );
buf1 gate1416( .a(N4599), .O(N4697) );
buf1 gate1417( .a(N4599), .O(N4700) );
inv1 gate( .a(N4629),.O(N4629_NOT) );
inv1 gate( .a(N4668),.O(N4668_NOT));
and2 gate( .a(N4629_NOT), .b(p553), .O(EX1381) );
and2 gate( .a(N4668_NOT), .b(EX1381), .O(EX1382) );
and2 gate( .a(N4629), .b(p554), .O(EX1383) );
and2 gate( .a(N4668_NOT), .b(EX1383), .O(EX1384) );
and2 gate( .a(N4629_NOT), .b(p555), .O(EX1385) );
and2 gate( .a(N4668), .b(EX1385), .O(EX1386) );
and2 gate( .a(N4629), .b(p556), .O(EX1387) );
and2 gate( .a(N4668), .b(EX1387), .O(EX1388) );
or2  gate( .a(EX1382), .b(EX1384), .O(EX1389) );
or2  gate( .a(EX1386), .b(EX1389), .O(EX1390) );
or2  gate( .a(EX1388), .b(EX1390), .O(N4704) );
nand2 gate1419( .a(N4139), .b(N4669), .O(N4705) );
inv1 gate1420( .a(N4656), .O(N4706) );
inv1 gate1421( .a(N4659), .O(N4707) );
inv1 gate( .a(N4435),.O(N4435_NOT) );
inv1 gate( .a(N4673),.O(N4673_NOT));
and2 gate( .a(N4435_NOT), .b(p557), .O(EX1391) );
and2 gate( .a(N4673_NOT), .b(EX1391), .O(EX1392) );
and2 gate( .a(N4435), .b(p558), .O(EX1393) );
and2 gate( .a(N4673_NOT), .b(EX1393), .O(EX1394) );
and2 gate( .a(N4435_NOT), .b(p559), .O(EX1395) );
and2 gate( .a(N4673), .b(EX1395), .O(EX1396) );
and2 gate( .a(N4435), .b(p560), .O(EX1397) );
and2 gate( .a(N4673), .b(EX1397), .O(EX1398) );
or2  gate( .a(EX1392), .b(EX1394), .O(EX1399) );
or2  gate( .a(EX1396), .b(EX1399), .O(EX1400) );
or2  gate( .a(EX1398), .b(EX1400), .O(N4708) );
nand2 gate1423( .a(N4675), .b(N4636), .O(N4711) );
inv1 gate( .a(N4493),.O(N4493_NOT) );
inv1 gate( .a(N4676),.O(N4676_NOT));
and2 gate( .a(N4493_NOT), .b(p561), .O(EX1401) );
and2 gate( .a(N4676_NOT), .b(EX1401), .O(EX1402) );
and2 gate( .a(N4493), .b(p562), .O(EX1403) );
and2 gate( .a(N4676_NOT), .b(EX1403), .O(EX1404) );
and2 gate( .a(N4493_NOT), .b(p563), .O(EX1405) );
and2 gate( .a(N4676), .b(EX1405), .O(EX1406) );
and2 gate( .a(N4493), .b(p564), .O(EX1407) );
and2 gate( .a(N4676), .b(EX1407), .O(EX1408) );
or2  gate( .a(EX1402), .b(EX1404), .O(EX1409) );
or2  gate( .a(EX1406), .b(EX1409), .O(EX1410) );
or2  gate( .a(EX1408), .b(EX1410), .O(N4716) );
nand2 gate1425( .a(N4678), .b(N4641), .O(N4717) );
nand2 gate1426( .a(N4679), .b(N4643), .O(N4721) );
buf1 gate1427( .a(N4644), .O(N4722) );
inv1 gate1428( .a(N4664), .O(N4726) );
or3 gate1429( .a(N4647), .b(N4650), .c(N4350), .O(N4727) );
nor3 gate1430( .a(N4647), .b(N4650), .c(N4350), .O(N4730) );
nand2 gate1431( .a(N4479), .b(N4687), .O(N4733) );
nand2 gate1432( .a(N4705), .b(N4670), .O(N4740) );
nand2 gate1433( .a(N4708), .b(N4674), .O(N4743) );
inv1 gate1434( .a(N4691), .O(N4747) );
nand2 gate1435( .a(N4691), .b(N4596), .O(N4748) );
inv1 gate1436( .a(N4694), .O(N4749) );
nand2 gate1437( .a(N4694), .b(N4597), .O(N4750) );
inv1 gate1438( .a(N4697), .O(N4753) );
nand2 gate1439( .a(N4697), .b(N4602), .O(N4754) );
inv1 gate1440( .a(N4700), .O(N4755) );
nand2 gate1441( .a(N4700), .b(N4603), .O(N4756) );
nand2 gate1442( .a(N4716), .b(N4677), .O(N4757) );
nand2 gate1443( .a(N4733), .b(N4688), .O(N4769) );
and2 gate1444( .a(N330), .b(N4704), .O(N4772) );
inv1 gate1445( .a(N4721), .O(N4775) );
inv1 gate1446( .a(N4730), .O(N4778) );
inv1 gate( .a(N4531),.O(N4531_NOT) );
inv1 gate( .a(N4747),.O(N4747_NOT));
and2 gate( .a(N4531_NOT), .b(p565), .O(EX1411) );
and2 gate( .a(N4747_NOT), .b(EX1411), .O(EX1412) );
and2 gate( .a(N4531), .b(p566), .O(EX1413) );
and2 gate( .a(N4747_NOT), .b(EX1413), .O(EX1414) );
and2 gate( .a(N4531_NOT), .b(p567), .O(EX1415) );
and2 gate( .a(N4747), .b(EX1415), .O(EX1416) );
and2 gate( .a(N4531), .b(p568), .O(EX1417) );
and2 gate( .a(N4747), .b(EX1417), .O(EX1418) );
or2  gate( .a(EX1412), .b(EX1414), .O(EX1419) );
or2  gate( .a(EX1416), .b(EX1419), .O(EX1420) );
or2  gate( .a(EX1418), .b(EX1420), .O(N4786) );
nand2 gate1448( .a(N4534), .b(N4749), .O(N4787) );
nand2 gate1449( .a(N4537), .b(N4753), .O(N4788) );
nand2 gate1450( .a(N4540), .b(N4755), .O(N4789) );
and2 gate1451( .a(N4711), .b(N2124), .O(N4794) );
inv1 gate( .a(N4711),.O(N4711_NOT) );
inv1 gate( .a(N2735),.O(N2735_NOT));
and2 gate( .a(N4711_NOT), .b(p569), .O(EX1421) );
and2 gate( .a(N2735_NOT), .b(EX1421), .O(EX1422) );
and2 gate( .a(N4711), .b(p570), .O(EX1423) );
and2 gate( .a(N2735_NOT), .b(EX1423), .O(EX1424) );
and2 gate( .a(N4711_NOT), .b(p571), .O(EX1425) );
and2 gate( .a(N2735), .b(EX1425), .O(EX1426) );
and2 gate( .a(N4711), .b(p572), .O(EX1427) );
and2 gate( .a(N2735), .b(EX1427), .O(EX1428) );
or2  gate( .a(EX1422), .b(EX1424), .O(EX1429) );
or2  gate( .a(EX1426), .b(EX1429), .O(EX1430) );
or2  gate( .a(EX1428), .b(EX1430), .O(N4797) );
and2 gate1453( .a(N4717), .b(N2127), .O(N4800) );
buf1 gate1454( .a(N4722), .O(N4805) );
inv1 gate( .a(N4717),.O(N4717_NOT) );
inv1 gate( .a(N4468),.O(N4468_NOT));
and2 gate( .a(N4717_NOT), .b(p573), .O(EX1431) );
and2 gate( .a(N4468_NOT), .b(EX1431), .O(EX1432) );
and2 gate( .a(N4717), .b(p574), .O(EX1433) );
and2 gate( .a(N4468_NOT), .b(EX1433), .O(EX1434) );
and2 gate( .a(N4717_NOT), .b(p575), .O(EX1435) );
and2 gate( .a(N4468), .b(EX1435), .O(EX1436) );
and2 gate( .a(N4717), .b(p576), .O(EX1437) );
and2 gate( .a(N4468), .b(EX1437), .O(EX1438) );
or2  gate( .a(EX1432), .b(EX1434), .O(EX1439) );
or2  gate( .a(EX1436), .b(EX1439), .O(EX1440) );
or2  gate( .a(EX1438), .b(EX1440), .O(N4808) );
buf1 gate1456( .a(N4727), .O(N4812) );
and2 gate1457( .a(N4727), .b(N4778), .O(N4815) );
inv1 gate1458( .a(N4769), .O(N4816) );
inv1 gate1459( .a(N4772), .O(N4817) );
inv1 gate( .a(N4786),.O(N4786_NOT) );
inv1 gate( .a(N4748),.O(N4748_NOT));
and2 gate( .a(N4786_NOT), .b(p577), .O(EX1441) );
and2 gate( .a(N4748_NOT), .b(EX1441), .O(EX1442) );
and2 gate( .a(N4786), .b(p578), .O(EX1443) );
and2 gate( .a(N4748_NOT), .b(EX1443), .O(EX1444) );
and2 gate( .a(N4786_NOT), .b(p579), .O(EX1445) );
and2 gate( .a(N4748), .b(EX1445), .O(EX1446) );
and2 gate( .a(N4786), .b(p580), .O(EX1447) );
and2 gate( .a(N4748), .b(EX1447), .O(EX1448) );
or2  gate( .a(EX1442), .b(EX1444), .O(EX1449) );
or2  gate( .a(EX1446), .b(EX1449), .O(EX1450) );
or2  gate( .a(EX1448), .b(EX1450), .O(N4818) );
nand2 gate1461( .a(N4787), .b(N4750), .O(N4822) );
nand2 gate1462( .a(N4788), .b(N4754), .O(N4823) );
nand2 gate1463( .a(N4789), .b(N4756), .O(N4826) );
nand2 gate1464( .a(N4775), .b(N4726), .O(N4829) );
inv1 gate1465( .a(N4775), .O(N4830) );
and2 gate1466( .a(N4743), .b(N2122), .O(N4831) );
and2 gate1467( .a(N4757), .b(N2126), .O(N4838) );
buf1 gate1468( .a(N4740), .O(N4844) );
buf1 gate1469( .a(N4740), .O(N4847) );
buf1 gate1470( .a(N4743), .O(N4850) );
buf1 gate1471( .a(N4757), .O(N4854) );
nand2 gate1472( .a(N4772), .b(N4816), .O(N4859) );
nand2 gate1473( .a(N4769), .b(N4817), .O(N4860) );
inv1 gate1474( .a(N4826), .O(N4868) );
inv1 gate1475( .a(N4805), .O(N4870) );
inv1 gate1476( .a(N4808), .O(N4872) );
nand2 gate1477( .a(N4664), .b(N4830), .O(N4873) );
or3 gate1478( .a(N4794), .b(N4797), .c(N4341), .O(N4876) );
nor3 gate1479( .a(N4794), .b(N4797), .c(N4341), .O(N4880) );
inv1 gate1480( .a(N4812), .O(N4885) );
inv1 gate1481( .a(N4822), .O(N4889) );
nand2 gate1482( .a(N4859), .b(N4860), .O(N4895) );
inv1 gate1483( .a(N4844), .O(N4896) );
nand2 gate1484( .a(N4844), .b(N4706), .O(N4897) );
inv1 gate1485( .a(N4847), .O(N4898) );
nand2 gate1486( .a(N4847), .b(N4707), .O(N4899) );
nor2 gate1487( .a(N4868), .b(N4564), .O(N4900) );
and4 gate1488( .a(N4717), .b(N4757), .c(N4823), .d(N4564), .O(N4901) );
inv1 gate1489( .a(N4850), .O(N4902) );
inv1 gate1490( .a(N4854), .O(N4904) );
inv1 gate( .a(N4854),.O(N4854_NOT) );
inv1 gate( .a(N4872),.O(N4872_NOT));
and2 gate( .a(N4854_NOT), .b(p581), .O(EX1451) );
and2 gate( .a(N4872_NOT), .b(EX1451), .O(EX1452) );
and2 gate( .a(N4854), .b(p582), .O(EX1453) );
and2 gate( .a(N4872_NOT), .b(EX1453), .O(EX1454) );
and2 gate( .a(N4854_NOT), .b(p583), .O(EX1455) );
and2 gate( .a(N4872), .b(EX1455), .O(EX1456) );
and2 gate( .a(N4854), .b(p584), .O(EX1457) );
and2 gate( .a(N4872), .b(EX1457), .O(EX1458) );
or2  gate( .a(EX1452), .b(EX1454), .O(EX1459) );
or2  gate( .a(EX1456), .b(EX1459), .O(EX1460) );
or2  gate( .a(EX1458), .b(EX1460), .O(N4905) );
nand2 gate1492( .a(N4873), .b(N4829), .O(N4906) );
and2 gate1493( .a(N4818), .b(N2123), .O(N4907) );
and2 gate1494( .a(N4823), .b(N2125), .O(N4913) );
and2 gate1495( .a(N4818), .b(N4644), .O(N4916) );
inv1 gate1496( .a(N4880), .O(N4920) );
inv1 gate( .a(N4895),.O(N4895_NOT) );
inv1 gate( .a(N2184),.O(N2184_NOT));
and2 gate( .a(N4895_NOT), .b(p585), .O(EX1461) );
and2 gate( .a(N2184_NOT), .b(EX1461), .O(EX1462) );
and2 gate( .a(N4895), .b(p586), .O(EX1463) );
and2 gate( .a(N2184_NOT), .b(EX1463), .O(EX1464) );
and2 gate( .a(N4895_NOT), .b(p587), .O(EX1465) );
and2 gate( .a(N2184), .b(EX1465), .O(EX1466) );
and2 gate( .a(N4895), .b(p588), .O(EX1467) );
and2 gate( .a(N2184), .b(EX1467), .O(EX1468) );
or2  gate( .a(EX1462), .b(EX1464), .O(EX1469) );
or2  gate( .a(EX1466), .b(EX1469), .O(EX1470) );
or2  gate( .a(EX1468), .b(EX1470), .O(N4921) );
nand2 gate1498( .a(N4656), .b(N4896), .O(N4924) );
nand2 gate1499( .a(N4659), .b(N4898), .O(N4925) );
or2 gate1500( .a(N4900), .b(N4901), .O(N4926) );
nand2 gate1501( .a(N4889), .b(N4870), .O(N4928) );
inv1 gate1502( .a(N4889), .O(N4929) );
nand2 gate1503( .a(N4808), .b(N4904), .O(N4930) );
inv1 gate1504( .a(N4906), .O(N4931) );
buf1 gate1505( .a(N4876), .O(N4937) );
buf1 gate1506( .a(N4876), .O(N4940) );
and2 gate1507( .a(N4876), .b(N4920), .O(N4944) );
nand2 gate1508( .a(N4924), .b(N4897), .O(N4946) );
nand2 gate1509( .a(N4925), .b(N4899), .O(N4949) );
nand2 gate1510( .a(N4916), .b(N4902), .O(N4950) );
inv1 gate1511( .a(N4916), .O(N4951) );
nand2 gate1512( .a(N4805), .b(N4929), .O(N4952) );
inv1 gate( .a(N4930),.O(N4930_NOT) );
inv1 gate( .a(N4905),.O(N4905_NOT));
and2 gate( .a(N4930_NOT), .b(p589), .O(EX1471) );
and2 gate( .a(N4905_NOT), .b(EX1471), .O(EX1472) );
and2 gate( .a(N4930), .b(p590), .O(EX1473) );
and2 gate( .a(N4905_NOT), .b(EX1473), .O(EX1474) );
and2 gate( .a(N4930_NOT), .b(p591), .O(EX1475) );
and2 gate( .a(N4905), .b(EX1475), .O(EX1476) );
and2 gate( .a(N4930), .b(p592), .O(EX1477) );
and2 gate( .a(N4905), .b(EX1477), .O(EX1478) );
or2  gate( .a(EX1472), .b(EX1474), .O(EX1479) );
or2  gate( .a(EX1476), .b(EX1479), .O(EX1480) );
or2  gate( .a(EX1478), .b(EX1480), .O(N4953) );
and2 gate1514( .a(N4926), .b(N2737), .O(N4954) );
and2 gate1515( .a(N4931), .b(N2741), .O(N4957) );
or3 gate1516( .a(N2764), .b(N2483), .c(N4921), .O(N4964) );
nor3 gate1517( .a(N2764), .b(N2483), .c(N4921), .O(N4965) );
inv1 gate1518( .a(N4949), .O(N4968) );
nand2 gate1519( .a(N4850), .b(N4951), .O(N4969) );
nand2 gate1520( .a(N4952), .b(N4928), .O(N4970) );
inv1 gate( .a(N4953),.O(N4953_NOT) );
inv1 gate( .a(N2739),.O(N2739_NOT));
and2 gate( .a(N4953_NOT), .b(p593), .O(EX1481) );
and2 gate( .a(N2739_NOT), .b(EX1481), .O(EX1482) );
and2 gate( .a(N4953), .b(p594), .O(EX1483) );
and2 gate( .a(N2739_NOT), .b(EX1483), .O(EX1484) );
and2 gate( .a(N4953_NOT), .b(p595), .O(EX1485) );
and2 gate( .a(N2739), .b(EX1485), .O(EX1486) );
and2 gate( .a(N4953), .b(p596), .O(EX1487) );
and2 gate( .a(N2739), .b(EX1487), .O(EX1488) );
or2  gate( .a(EX1482), .b(EX1484), .O(EX1489) );
or2  gate( .a(EX1486), .b(EX1489), .O(EX1490) );
or2  gate( .a(EX1488), .b(EX1490), .O(N4973) );
inv1 gate1522( .a(N4937), .O(N4978) );
inv1 gate1523( .a(N4940), .O(N4979) );
inv1 gate1524( .a(N4965), .O(N4980) );
nor2 gate1525( .a(N4968), .b(N4722), .O(N4981) );
and4 gate1526( .a(N4818), .b(N4743), .c(N4946), .d(N4722), .O(N4982) );
inv1 gate( .a(N4950),.O(N4950_NOT) );
inv1 gate( .a(N4969),.O(N4969_NOT));
and2 gate( .a(N4950_NOT), .b(p597), .O(EX1491) );
and2 gate( .a(N4969_NOT), .b(EX1491), .O(EX1492) );
and2 gate( .a(N4950), .b(p598), .O(EX1493) );
and2 gate( .a(N4969_NOT), .b(EX1493), .O(EX1494) );
and2 gate( .a(N4950_NOT), .b(p599), .O(EX1495) );
and2 gate( .a(N4969), .b(EX1495), .O(EX1496) );
and2 gate( .a(N4950), .b(p600), .O(EX1497) );
and2 gate( .a(N4969), .b(EX1497), .O(EX1498) );
or2  gate( .a(EX1492), .b(EX1494), .O(EX1499) );
or2  gate( .a(EX1496), .b(EX1499), .O(EX1500) );
or2  gate( .a(EX1498), .b(EX1500), .O(N4983) );
inv1 gate1528( .a(N4970), .O(N4984) );
and2 gate1529( .a(N4946), .b(N2121), .O(N4985) );
or3 gate1530( .a(N4913), .b(N4954), .c(N4344), .O(N4988) );
nor3 gate1531( .a(N4913), .b(N4954), .c(N4344), .O(N4991) );
or3 gate1532( .a(N4800), .b(N4957), .c(N4347), .O(N4996) );
nor3 gate1533( .a(N4800), .b(N4957), .c(N4347), .O(N4999) );
and2 gate1534( .a(N4964), .b(N4980), .O(N5002) );
inv1 gate( .a(N4981),.O(N4981_NOT) );
inv1 gate( .a(N4982),.O(N4982_NOT));
and2 gate( .a(N4981_NOT), .b(p601), .O(EX1501) );
and2 gate( .a(N4982_NOT), .b(EX1501), .O(EX1502) );
and2 gate( .a(N4981), .b(p602), .O(EX1503) );
and2 gate( .a(N4982_NOT), .b(EX1503), .O(EX1504) );
and2 gate( .a(N4981_NOT), .b(p603), .O(EX1505) );
and2 gate( .a(N4982), .b(EX1505), .O(EX1506) );
and2 gate( .a(N4981), .b(p604), .O(EX1507) );
and2 gate( .a(N4982), .b(EX1507), .O(EX1508) );
or2  gate( .a(EX1502), .b(EX1504), .O(EX1509) );
or2  gate( .a(EX1506), .b(EX1509), .O(EX1510) );
or2  gate( .a(EX1508), .b(EX1510), .O(N5007) );
and2 gate1536( .a(N4983), .b(N2731), .O(N5010) );
and2 gate1537( .a(N4984), .b(N2733), .O(N5013) );
or3 gate1538( .a(N4838), .b(N4973), .c(N4475), .O(N5018) );
nor3 gate1539( .a(N4838), .b(N4973), .c(N4475), .O(N5021) );
inv1 gate1540( .a(N4991), .O(N5026) );
inv1 gate1541( .a(N4999), .O(N5029) );
inv1 gate( .a(N5007),.O(N5007_NOT) );
inv1 gate( .a(N2729),.O(N2729_NOT));
and2 gate( .a(N5007_NOT), .b(p605), .O(EX1511) );
and2 gate( .a(N2729_NOT), .b(EX1511), .O(EX1512) );
and2 gate( .a(N5007), .b(p606), .O(EX1513) );
and2 gate( .a(N2729_NOT), .b(EX1513), .O(EX1514) );
and2 gate( .a(N5007_NOT), .b(p607), .O(EX1515) );
and2 gate( .a(N2729), .b(EX1515), .O(EX1516) );
and2 gate( .a(N5007), .b(p608), .O(EX1517) );
and2 gate( .a(N2729), .b(EX1517), .O(EX1518) );
or2  gate( .a(EX1512), .b(EX1514), .O(EX1519) );
or2  gate( .a(EX1516), .b(EX1519), .O(EX1520) );
or2  gate( .a(EX1518), .b(EX1520), .O(N5030) );
buf1 gate1543( .a(N4996), .O(N5039) );
buf1 gate1544( .a(N4988), .O(N5042) );
and2 gate1545( .a(N4988), .b(N5026), .O(N5045) );
inv1 gate1546( .a(N5021), .O(N5046) );
and2 gate1547( .a(N4996), .b(N5029), .O(N5047) );
or3 gate1548( .a(N4831), .b(N5010), .c(N4472), .O(N5050) );
nor3 gate1549( .a(N4831), .b(N5010), .c(N4472), .O(N5055) );
or3 gate1550( .a(N4907), .b(N5013), .c(N4338), .O(N5058) );
nor3 gate1551( .a(N4907), .b(N5013), .c(N4338), .O(N5061) );
and4 gate1552( .a(N4730), .b(N4999), .c(N5021), .d(N4991), .O(N5066) );
buf1 gate1553( .a(N5018), .O(N5070) );
and2 gate1554( .a(N5018), .b(N5046), .O(N5078) );
or3 gate1555( .a(N4985), .b(N5030), .c(N4335), .O(N5080) );
nor3 gate1556( .a(N4985), .b(N5030), .c(N4335), .O(N5085) );
nand2 gate1557( .a(N5039), .b(N4885), .O(N5094) );
inv1 gate1558( .a(N5039), .O(N5095) );
inv1 gate1559( .a(N5042), .O(N5097) );
inv1 gate( .a(N5050),.O(N5050_NOT) );
inv1 gate( .a(N5050),.O(N5050_NOT));
and2 gate( .a(N5050_NOT), .b(p609), .O(EX1521) );
and2 gate( .a(N5050_NOT), .b(EX1521), .O(EX1522) );
and2 gate( .a(N5050), .b(p610), .O(EX1523) );
and2 gate( .a(N5050_NOT), .b(EX1523), .O(EX1524) );
and2 gate( .a(N5050_NOT), .b(p611), .O(EX1525) );
and2 gate( .a(N5050), .b(EX1525), .O(EX1526) );
and2 gate( .a(N5050), .b(p612), .O(EX1527) );
and2 gate( .a(N5050), .b(EX1527), .O(EX1528) );
or2  gate( .a(EX1522), .b(EX1524), .O(EX1529) );
or2  gate( .a(EX1526), .b(EX1529), .O(EX1530) );
or2  gate( .a(EX1528), .b(EX1530), .O(N5102) );
inv1 gate1561( .a(N5061), .O(N5103) );
nand2 gate1562( .a(N4812), .b(N5095), .O(N5108) );
inv1 gate1563( .a(N5070), .O(N5109) );
nand2 gate1564( .a(N5070), .b(N5097), .O(N5110) );
buf1 gate1565( .a(N5058), .O(N5111) );
and2 gate1566( .a(N5050), .b(N1461), .O(N5114) );
buf1 gate1567( .a(N5050), .O(N5117) );
and2 gate1568( .a(N5080), .b(N5080), .O(N5120) );
and2 gate1569( .a(N5058), .b(N5103), .O(N5121) );
nand2 gate1570( .a(N5094), .b(N5108), .O(N5122) );
nand2 gate1571( .a(N5042), .b(N5109), .O(N5125) );
inv1 gate( .a(N1461),.O(N1461_NOT) );
inv1 gate( .a(N5080),.O(N5080_NOT));
and2 gate( .a(N1461_NOT), .b(p613), .O(EX1531) );
and2 gate( .a(N5080_NOT), .b(EX1531), .O(EX1532) );
and2 gate( .a(N1461), .b(p614), .O(EX1533) );
and2 gate( .a(N5080_NOT), .b(EX1533), .O(EX1534) );
and2 gate( .a(N1461_NOT), .b(p615), .O(EX1535) );
and2 gate( .a(N5080), .b(EX1535), .O(EX1536) );
and2 gate( .a(N1461), .b(p616), .O(EX1537) );
and2 gate( .a(N5080), .b(EX1537), .O(EX1538) );
or2  gate( .a(EX1532), .b(EX1534), .O(EX1539) );
or2  gate( .a(EX1536), .b(EX1539), .O(EX1540) );
or2  gate( .a(EX1538), .b(EX1540), .O(N5128) );
and4 gate1573( .a(N4880), .b(N5061), .c(N5055), .d(N5085), .O(N5133) );
and3 gate1574( .a(N5055), .b(N5085), .c(N1464), .O(N5136) );
buf1 gate1575( .a(N5080), .O(N5139) );
nand2 gate1576( .a(N5125), .b(N5110), .O(N5145) );
buf1 gate1577( .a(N5111), .O(N5151) );
buf1 gate1578( .a(N5111), .O(N5154) );
inv1 gate1579( .a(N5117), .O(N5159) );
buf1 gate1580( .a(N5114), .O(N5160) );
buf1 gate1581( .a(N5114), .O(N5163) );
and2 gate1582( .a(N5066), .b(N5133), .O(N5166) );
and2 gate1583( .a(N5066), .b(N5133), .O(N5173) );
buf1 gate1584( .a(N5122), .O(N5174) );
buf1 gate1585( .a(N5122), .O(N5177) );
inv1 gate1586( .a(N5139), .O(N5182) );
nand2 gate1587( .a(N5139), .b(N5159), .O(N5183) );
buf1 gate1588( .a(N5128), .O(N5184) );
buf1 gate1589( .a(N5128), .O(N5188) );
inv1 gate1590( .a(N5166), .O(N5192) );
nor2 gate1591( .a(N5136), .b(N5173), .O(N5193) );
nand2 gate1592( .a(N5151), .b(N4978), .O(N5196) );
inv1 gate1593( .a(N5151), .O(N5197) );
nand2 gate1594( .a(N5154), .b(N4979), .O(N5198) );
inv1 gate1595( .a(N5154), .O(N5199) );
inv1 gate1596( .a(N5160), .O(N5201) );
inv1 gate1597( .a(N5163), .O(N5203) );
buf1 gate1598( .a(N5145), .O(N5205) );
buf1 gate1599( .a(N5145), .O(N5209) );
nand2 gate1600( .a(N5117), .b(N5182), .O(N5212) );
inv1 gate( .a(N213),.O(N213_NOT) );
inv1 gate( .a(N5193),.O(N5193_NOT));
and2 gate( .a(N213_NOT), .b(p617), .O(EX1541) );
and2 gate( .a(N5193_NOT), .b(EX1541), .O(EX1542) );
and2 gate( .a(N213), .b(p618), .O(EX1543) );
and2 gate( .a(N5193_NOT), .b(EX1543), .O(EX1544) );
and2 gate( .a(N213_NOT), .b(p619), .O(EX1545) );
and2 gate( .a(N5193), .b(EX1545), .O(EX1546) );
and2 gate( .a(N213), .b(p620), .O(EX1547) );
and2 gate( .a(N5193), .b(EX1547), .O(EX1548) );
or2  gate( .a(EX1542), .b(EX1544), .O(EX1549) );
or2  gate( .a(EX1546), .b(EX1549), .O(EX1550) );
or2  gate( .a(EX1548), .b(EX1550), .O(N5215) );
inv1 gate1602( .a(N5174), .O(N5217) );
inv1 gate1603( .a(N5177), .O(N5219) );
inv1 gate( .a(N4937),.O(N4937_NOT) );
inv1 gate( .a(N5197),.O(N5197_NOT));
and2 gate( .a(N4937_NOT), .b(p621), .O(EX1551) );
and2 gate( .a(N5197_NOT), .b(EX1551), .O(EX1552) );
and2 gate( .a(N4937), .b(p622), .O(EX1553) );
and2 gate( .a(N5197_NOT), .b(EX1553), .O(EX1554) );
and2 gate( .a(N4937_NOT), .b(p623), .O(EX1555) );
and2 gate( .a(N5197), .b(EX1555), .O(EX1556) );
and2 gate( .a(N4937), .b(p624), .O(EX1557) );
and2 gate( .a(N5197), .b(EX1557), .O(EX1558) );
or2  gate( .a(EX1552), .b(EX1554), .O(EX1559) );
or2  gate( .a(EX1556), .b(EX1559), .O(EX1560) );
or2  gate( .a(EX1558), .b(EX1560), .O(N5220) );
nand2 gate1605( .a(N4940), .b(N5199), .O(N5221) );
inv1 gate1606( .a(N5184), .O(N5222) );
nand2 gate1607( .a(N5184), .b(N5201), .O(N5223) );
nand2 gate1608( .a(N5188), .b(N5203), .O(N5224) );
inv1 gate1609( .a(N5188), .O(N5225) );
nand2 gate1610( .a(N5183), .b(N5212), .O(N5228) );
inv1 gate1611( .a(N5215), .O(N5231) );
inv1 gate( .a(N5205),.O(N5205_NOT) );
inv1 gate( .a(N5217),.O(N5217_NOT));
and2 gate( .a(N5205_NOT), .b(p625), .O(EX1561) );
and2 gate( .a(N5217_NOT), .b(EX1561), .O(EX1562) );
and2 gate( .a(N5205), .b(p626), .O(EX1563) );
and2 gate( .a(N5217_NOT), .b(EX1563), .O(EX1564) );
and2 gate( .a(N5205_NOT), .b(p627), .O(EX1565) );
and2 gate( .a(N5217), .b(EX1565), .O(EX1566) );
and2 gate( .a(N5205), .b(p628), .O(EX1567) );
and2 gate( .a(N5217), .b(EX1567), .O(EX1568) );
or2  gate( .a(EX1562), .b(EX1564), .O(EX1569) );
or2  gate( .a(EX1566), .b(EX1569), .O(EX1570) );
or2  gate( .a(EX1568), .b(EX1570), .O(N5232) );
inv1 gate1613( .a(N5205), .O(N5233) );
nand2 gate1614( .a(N5209), .b(N5219), .O(N5234) );
inv1 gate1615( .a(N5209), .O(N5235) );
nand2 gate1616( .a(N5196), .b(N5220), .O(N5236) );
inv1 gate( .a(N5198),.O(N5198_NOT) );
inv1 gate( .a(N5221),.O(N5221_NOT));
and2 gate( .a(N5198_NOT), .b(p629), .O(EX1571) );
and2 gate( .a(N5221_NOT), .b(EX1571), .O(EX1572) );
and2 gate( .a(N5198), .b(p630), .O(EX1573) );
and2 gate( .a(N5221_NOT), .b(EX1573), .O(EX1574) );
and2 gate( .a(N5198_NOT), .b(p631), .O(EX1575) );
and2 gate( .a(N5221), .b(EX1575), .O(EX1576) );
and2 gate( .a(N5198), .b(p632), .O(EX1577) );
and2 gate( .a(N5221), .b(EX1577), .O(EX1578) );
or2  gate( .a(EX1572), .b(EX1574), .O(EX1579) );
or2  gate( .a(EX1576), .b(EX1579), .O(EX1580) );
or2  gate( .a(EX1578), .b(EX1580), .O(N5240) );
nand2 gate1618( .a(N5160), .b(N5222), .O(N5242) );
nand2 gate1619( .a(N5163), .b(N5225), .O(N5243) );
nand2 gate1620( .a(N5174), .b(N5233), .O(N5245) );
nand2 gate1621( .a(N5177), .b(N5235), .O(N5246) );
inv1 gate1622( .a(N5240), .O(N5250) );
inv1 gate1623( .a(N5228), .O(N5253) );
nand2 gate1624( .a(N5242), .b(N5223), .O(N5254) );
nand2 gate1625( .a(N5243), .b(N5224), .O(N5257) );
inv1 gate( .a(N5232),.O(N5232_NOT) );
inv1 gate( .a(N5245),.O(N5245_NOT));
and2 gate( .a(N5232_NOT), .b(p633), .O(EX1581) );
and2 gate( .a(N5245_NOT), .b(EX1581), .O(EX1582) );
and2 gate( .a(N5232), .b(p634), .O(EX1583) );
and2 gate( .a(N5245_NOT), .b(EX1583), .O(EX1584) );
and2 gate( .a(N5232_NOT), .b(p635), .O(EX1585) );
and2 gate( .a(N5245), .b(EX1585), .O(EX1586) );
and2 gate( .a(N5232), .b(p636), .O(EX1587) );
and2 gate( .a(N5245), .b(EX1587), .O(EX1588) );
or2  gate( .a(EX1582), .b(EX1584), .O(EX1589) );
or2  gate( .a(EX1586), .b(EX1589), .O(EX1590) );
or2  gate( .a(EX1588), .b(EX1590), .O(N5258) );
nand2 gate1627( .a(N5234), .b(N5246), .O(N5261) );
inv1 gate1628( .a(N5257), .O(N5266) );
buf1 gate1629( .a(N5236), .O(N5269) );
and3 gate1630( .a(N5236), .b(N5254), .c(N2307), .O(N5277) );
and3 gate1631( .a(N5250), .b(N5254), .c(N2310), .O(N5278) );
inv1 gate1632( .a(N5261), .O(N5279) );
inv1 gate1633( .a(N5269), .O(N5283) );
nand2 gate1634( .a(N5269), .b(N5253), .O(N5284) );
and3 gate1635( .a(N5236), .b(N5266), .c(N2310), .O(N5285) );
and3 gate1636( .a(N5250), .b(N5266), .c(N2307), .O(N5286) );
buf1 gate1637( .a(N5258), .O(N5289) );
buf1 gate1638( .a(N5258), .O(N5292) );
nand2 gate1639( .a(N5228), .b(N5283), .O(N5295) );
or4 gate1640( .a(N5277), .b(N5285), .c(N5278), .d(N5286), .O(N5298) );
buf1 gate1641( .a(N5279), .O(N5303) );
buf1 gate1642( .a(N5279), .O(N5306) );
inv1 gate( .a(N5295),.O(N5295_NOT) );
inv1 gate( .a(N5284),.O(N5284_NOT));
and2 gate( .a(N5295_NOT), .b(p637), .O(EX1591) );
and2 gate( .a(N5284_NOT), .b(EX1591), .O(EX1592) );
and2 gate( .a(N5295), .b(p638), .O(EX1593) );
and2 gate( .a(N5284_NOT), .b(EX1593), .O(EX1594) );
and2 gate( .a(N5295_NOT), .b(p639), .O(EX1595) );
and2 gate( .a(N5284), .b(EX1595), .O(EX1596) );
and2 gate( .a(N5295), .b(p640), .O(EX1597) );
and2 gate( .a(N5284), .b(EX1597), .O(EX1598) );
or2  gate( .a(EX1592), .b(EX1594), .O(EX1599) );
or2  gate( .a(EX1596), .b(EX1599), .O(EX1600) );
or2  gate( .a(EX1598), .b(EX1600), .O(N5309) );
inv1 gate1644( .a(N5292), .O(N5312) );
inv1 gate1645( .a(N5289), .O(N5313) );
inv1 gate1646( .a(N5306), .O(N5322) );
inv1 gate1647( .a(N5303), .O(N5323) );
buf1 gate1648( .a(N5298), .O(N5324) );
buf1 gate1649( .a(N5298), .O(N5327) );
buf1 gate1650( .a(N5309), .O(N5332) );
buf1 gate1651( .a(N5309), .O(N5335) );
inv1 gate( .a(N5324),.O(N5324_NOT) );
inv1 gate( .a(N5323),.O(N5323_NOT));
and2 gate( .a(N5324_NOT), .b(p641), .O(EX1601) );
and2 gate( .a(N5323_NOT), .b(EX1601), .O(EX1602) );
and2 gate( .a(N5324), .b(p642), .O(EX1603) );
and2 gate( .a(N5323_NOT), .b(EX1603), .O(EX1604) );
and2 gate( .a(N5324_NOT), .b(p643), .O(EX1605) );
and2 gate( .a(N5323), .b(EX1605), .O(EX1606) );
and2 gate( .a(N5324), .b(p644), .O(EX1607) );
and2 gate( .a(N5323), .b(EX1607), .O(EX1608) );
or2  gate( .a(EX1602), .b(EX1604), .O(EX1609) );
or2  gate( .a(EX1606), .b(EX1609), .O(EX1610) );
or2  gate( .a(EX1608), .b(EX1610), .O(N5340) );
inv1 gate( .a(N5327),.O(N5327_NOT) );
inv1 gate( .a(N5322),.O(N5322_NOT));
and2 gate( .a(N5327_NOT), .b(p645), .O(EX1611) );
and2 gate( .a(N5322_NOT), .b(EX1611), .O(EX1612) );
and2 gate( .a(N5327), .b(p646), .O(EX1613) );
and2 gate( .a(N5322_NOT), .b(EX1613), .O(EX1614) );
and2 gate( .a(N5327_NOT), .b(p647), .O(EX1615) );
and2 gate( .a(N5322), .b(EX1615), .O(EX1616) );
and2 gate( .a(N5327), .b(p648), .O(EX1617) );
and2 gate( .a(N5322), .b(EX1617), .O(EX1618) );
or2  gate( .a(EX1612), .b(EX1614), .O(EX1619) );
or2  gate( .a(EX1616), .b(EX1619), .O(EX1620) );
or2  gate( .a(EX1618), .b(EX1620), .O(N5341) );
inv1 gate1654( .a(N5327), .O(N5344) );
inv1 gate1655( .a(N5324), .O(N5345) );
nand2 gate1656( .a(N5332), .b(N5313), .O(N5348) );
nand2 gate1657( .a(N5335), .b(N5312), .O(N5349) );
nand2 gate1658( .a(N5303), .b(N5345), .O(N5350) );
inv1 gate( .a(N5306),.O(N5306_NOT) );
inv1 gate( .a(N5344),.O(N5344_NOT));
and2 gate( .a(N5306_NOT), .b(p649), .O(EX1621) );
and2 gate( .a(N5344_NOT), .b(EX1621), .O(EX1622) );
and2 gate( .a(N5306), .b(p650), .O(EX1623) );
and2 gate( .a(N5344_NOT), .b(EX1623), .O(EX1624) );
and2 gate( .a(N5306_NOT), .b(p651), .O(EX1625) );
and2 gate( .a(N5344), .b(EX1625), .O(EX1626) );
and2 gate( .a(N5306), .b(p652), .O(EX1627) );
and2 gate( .a(N5344), .b(EX1627), .O(EX1628) );
or2  gate( .a(EX1622), .b(EX1624), .O(EX1629) );
or2  gate( .a(EX1626), .b(EX1629), .O(EX1630) );
or2  gate( .a(EX1628), .b(EX1630), .O(N5351) );
inv1 gate1660( .a(N5335), .O(N5352) );
inv1 gate1661( .a(N5332), .O(N5353) );
nand2 gate1662( .a(N5289), .b(N5353), .O(N5354) );
nand2 gate1663( .a(N5292), .b(N5352), .O(N5355) );
nand2 gate1664( .a(N5350), .b(N5340), .O(N5356) );
nand2 gate1665( .a(N5351), .b(N5341), .O(N5357) );
nand2 gate1666( .a(N5348), .b(N5354), .O(N5358) );
inv1 gate( .a(N5349),.O(N5349_NOT) );
inv1 gate( .a(N5355),.O(N5355_NOT));
and2 gate( .a(N5349_NOT), .b(p653), .O(EX1631) );
and2 gate( .a(N5355_NOT), .b(EX1631), .O(EX1632) );
and2 gate( .a(N5349), .b(p654), .O(EX1633) );
and2 gate( .a(N5355_NOT), .b(EX1633), .O(EX1634) );
and2 gate( .a(N5349_NOT), .b(p655), .O(EX1635) );
and2 gate( .a(N5355), .b(EX1635), .O(EX1636) );
and2 gate( .a(N5349), .b(p656), .O(EX1637) );
and2 gate( .a(N5355), .b(EX1637), .O(EX1638) );
or2  gate( .a(EX1632), .b(EX1634), .O(EX1639) );
or2  gate( .a(EX1636), .b(EX1639), .O(EX1640) );
or2  gate( .a(EX1638), .b(EX1640), .O(N5359) );
and2 gate1668( .a(N5356), .b(N5357), .O(N5360) );
nand2 gate1669( .a(N5358), .b(N5359), .O(N5361) );

xor2 gate( .a(X_1), .b(N50_new), .O(N50) );
xor2 gate( .a(X_2), .b(N58_new), .O(N58) );
xor2 gate( .a(X_3), .b(N68_new), .O(N68) );
xor2 gate( .a(X_4), .b(N77_new), .O(N77) );
xor2 gate( .a(X_5), .b(N87_new), .O(N87) );
xor2 gate( .a(X_6), .b(N97_new), .O(N97) );
xor2 gate( .a(X_7), .b(N107_new), .O(N107) );
xor2 gate( .a(X_8), .b(N116_new), .O(N116) );
xor2 gate( .a(X_9), .b(N257_new), .O(N257) );
xor2 gate( .a(X_10), .b(N264_new), .O(N264) );
xor2 gate( .a(X_11), .b(N1_new), .O(N1) );
xor2 gate( .a(X_12), .b(N13_new), .O(N13) );
xor2 gate( .a(X_13), .b(N20_new), .O(N20) );
xor2 gate( .a(X_14), .b(N33_new), .O(N33) );
xor2 gate( .a(X_15), .b(N41_new), .O(N41) );
xor2 gate( .a(X_16), .b(N45_new), .O(N45) );
xor2 gate( .a(X_17), .b(N190_new), .O(N190) );
xor2 gate( .a(X_18), .b(N200_new), .O(N200) );
xor2 gate( .a(X_19), .b(N179_new), .O(N179) );
xor2 gate( .a(X_20), .b(N349_new), .O(N349) );
xor2 gate( .a(X_21), .b(N213_new), .O(N213) );
xor2 gate( .a(X_22), .b(N343_new), .O(N343) );
xor2 gate( .a(X_23), .b(N226_new), .O(N226) );
xor2 gate( .a(X_24), .b(N232_new), .O(N232) );
xor2 gate( .a(X_25), .b(N238_new), .O(N238) );
xor2 gate( .a(X_26), .b(N244_new), .O(N244) );
xor2 gate( .a(X_27), .b(N250_new), .O(N250) );
xor2 gate( .a(X_28), .b(N270_new), .O(N270) );
xor2 gate( .a(X_29), .b(N330_new), .O(N330) );
xor2 gate( .a(X_30), .b(N169_new), .O(N169) );
xor2 gate( .a(X_31), .b(N222_new), .O(N222) );
xor2 gate( .a(X_32), .b(N223_new), .O(N223) );
xor2 gate( .a(X_33), .b(N1713), .O(N1713_new) );
xor2 gate( .a(X_34), .b(N150_new), .O(N150) );
xor2 gate( .a(X_35), .b(N159_new), .O(N159) );
xor2 gate( .a(X_36), .b(N283_new), .O(N283) );
xor2 gate( .a(X_37), .b(N1947), .O(N1947_new) );
xor2 gate( .a(X_38), .b(N294_new), .O(N294) );
xor2 gate( .a(X_39), .b(N303_new), .O(N303) );
xor2 gate( .a(X_40), .b(N350_new), .O(N350) );
xor2 gate( .a(X_41), .b(N274_new), .O(N274) );
xor2 gate( .a(X_42), .b(N3195), .O(N3195_new) );
xor2 gate( .a(X_43), .b(N124_new), .O(N124) );
xor2 gate( .a(X_44), .b(N143_new), .O(N143) );
xor2 gate( .a(X_45), .b(N137_new), .O(N137) );
xor2 gate( .a(X_46), .b(N132_new), .O(N132) );
xor2 gate( .a(X_47), .b(N128_new), .O(N128) );
xor2 gate( .a(X_48), .b(N125_new), .O(N125) );
xor2 gate( .a(X_49), .b(N311_new), .O(N311) );
xor2 gate( .a(X_50), .b(N317_new), .O(N317) );
xor2 gate( .a(X_51), .b(N322_new), .O(N322) );
xor2 gate( .a(X_52), .b(N326_new), .O(N326) );
xor2 gate( .a(X_53), .b(N329_new), .O(N329) );
xor2 gate( .a(X_54), .b(N3833), .O(N3833_new) );
xor2 gate( .a(X_55), .b(N3987), .O(N3987_new) );
xor2 gate( .a(X_56), .b(N4028), .O(N4028_new) );
xor2 gate( .a(X_57), .b(N4145), .O(N4145_new) );
xor2 gate( .a(X_58), .b(N4589), .O(N4589_new) );
xor2 gate( .a(X_59), .b(N4667), .O(N4667_new) );
xor2 gate( .a(X_60), .b(N4815), .O(N4815_new) );
xor2 gate( .a(X_61), .b(N4944), .O(N4944_new) );
xor2 gate( .a(X_62), .b(N5002), .O(N5002_new) );
xor2 gate( .a(X_63), .b(N5045), .O(N5045_new) );
xor2 gate( .a(X_64), .b(N5047), .O(N5047_new) );
xor2 gate( .a(X_65), .b(N5078), .O(N5078_new) );
xor2 gate( .a(X_66), .b(N5102), .O(N5102_new) );
xor2 gate( .a(X_67), .b(N5120), .O(N5120_new) );
xor2 gate( .a(X_68), .b(N5121), .O(N5121_new) );
xor2 gate( .a(X_69), .b(N5192), .O(N5192_new) );
xor2 gate( .a(X_70), .b(N5231), .O(N5231_new) );
xor2 gate( .a(X_71), .b(N5360), .O(N5360_new) );
xor2 gate( .a(X_72), .b(N5361), .O(N5361_new) );
endmodule