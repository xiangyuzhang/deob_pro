module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,             N753,N754,N755);


input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117_new,
      N121,N125,N129,N130,N131,N132,N133,N134,N135_new,N136,
      N137;

input p1,p2,p3,p4,X_1,X_2,X_3;


output N724,N725,N726,N727,N728,N729,N730,N731,N732_new,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;


wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,
     N288_NOT,N289_NOT,EX1,EX2,EX3,EX4,EX5,EX6,EX7,EX8,EX9,EX10,N135,N117,N732;

xor2 gate1( .a(N1), .b(N5), .O(N250) );
xor2 gate2( .a(N9), .b(N13), .O(N251) );
xor2 gate3( .a(N17), .b(N21), .O(N252) );
xor2 gate4( .a(N25), .b(N29), .O(N253) );
xor2 gate5( .a(N33), .b(N37), .O(N254) );
xor2 gate6( .a(N41), .b(N45), .O(N255) );
xor2 gate7( .a(N49), .b(N53), .O(N256) );
xor2 gate8( .a(N57), .b(N61), .O(N257) );
xor2 gate9( .a(N65), .b(N69), .O(N258) );
xor2 gate10( .a(N73), .b(N77), .O(N259) );
xor2 gate11( .a(N81), .b(N85), .O(N260) );
xor2 gate12( .a(N89), .b(N93), .O(N261) );
xor2 gate13( .a(N97), .b(N101), .O(N262) );
xor2 gate14( .a(N105), .b(N109), .O(N263) );
xor2 gate15( .a(N113), .b(N117), .O(N264) );
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );
xor2 gate26( .a(N33), .b(N49), .O(N275) );
xor2 gate27( .a(N5), .b(N21), .O(N276) );
xor2 gate28( .a(N37), .b(N53), .O(N277) );
xor2 gate29( .a(N9), .b(N25), .O(N278) );
xor2 gate30( .a(N41), .b(N57), .O(N279) );
xor2 gate31( .a(N13), .b(N29), .O(N280) );
xor2 gate32( .a(N45), .b(N61), .O(N281) );
xor2 gate33( .a(N65), .b(N81), .O(N282) );
xor2 gate34( .a(N97), .b(N113), .O(N283) );
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );
xor2 gate37( .a(N73), .b(N89), .O(N286) );
xor2 gate38( .a(N105), .b(N121), .O(N287) );
xor2 gate39( .a(N77), .b(N93), .O(N288) );
xor2 gate40( .a(N109), .b(N125), .O(N289) );
xor2 gate41( .a(N250), .b(N251), .O(N290) );
xor2 gate42( .a(N252), .b(N253), .O(N293) );
xor2 gate43( .a(N254), .b(N255), .O(N296) );
xor2 gate44( .a(N256), .b(N257), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );
xor2 gate46( .a(N260), .b(N261), .O(N305) );
xor2 gate47( .a(N262), .b(N263), .O(N308) );
xor2 gate48( .a(N264), .b(N265), .O(N311) );
xor2 gate49( .a(N274), .b(N275), .O(N314) );
xor2 gate50( .a(N276), .b(N277), .O(N315) );
xor2 gate51( .a(N278), .b(N279), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );
xor2 gate55( .a(N286), .b(N287), .O(N320) );
inv1 gate( .a(N288),.O(N288_NOT) );
inv1 gate( .a(N289),.O(N289_NOT));
and2 gate( .a(N288_NOT), .b(p1), .O(EX1) );
and2 gate( .a(N289_NOT), .b(EX1), .O(EX2) );
and2 gate( .a(N288), .b(p2), .O(EX3) );
and2 gate( .a(N289_NOT), .b(EX3), .O(EX4) );
and2 gate( .a(N288_NOT), .b(p3), .O(EX5) );
and2 gate( .a(N289), .b(EX5), .O(EX6) );
and2 gate( .a(N288), .b(p4), .O(EX7) );
and2 gate( .a(N289), .b(EX7), .O(EX8) );
or2  gate( .a(EX2), .b(EX4), .O(EX9) );
or2  gate( .a(EX6), .b(EX9), .O(EX10) );
or2  gate( .a(EX8), .b(EX10), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );
xor2 gate58( .a(N296), .b(N299), .O(N339) );
xor2 gate59( .a(N290), .b(N296), .O(N340) );
xor2 gate60( .a(N293), .b(N299), .O(N341) );
xor2 gate61( .a(N302), .b(N305), .O(N342) );
xor2 gate62( .a(N308), .b(N311), .O(N343) );
xor2 gate63( .a(N302), .b(N308), .O(N344) );
xor2 gate64( .a(N305), .b(N311), .O(N345) );
xor2 gate65( .a(N266), .b(N342), .O(N346) );
xor2 gate66( .a(N267), .b(N343), .O(N347) );
xor2 gate67( .a(N268), .b(N344), .O(N348) );
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );
xor2 gate70( .a(N271), .b(N339), .O(N351) );
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );
xor2 gate74( .a(N315), .b(N347), .O(N367) );
xor2 gate75( .a(N316), .b(N348), .O(N380) );
xor2 gate76( .a(N317), .b(N349), .O(N393) );
xor2 gate77( .a(N318), .b(N350), .O(N406) );
xor2 gate78( .a(N319), .b(N351), .O(N419) );
xor2 gate79( .a(N320), .b(N352), .O(N432) );
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );
xor2 gate172( .a(N5), .b(N693), .O(N725) );
xor2 gate173( .a(N9), .b(N694), .O(N726) );
xor2 gate174( .a(N13), .b(N695), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );
xor2 gate176( .a(N21), .b(N697), .O(N729) );
xor2 gate177( .a(N25), .b(N698), .O(N730) );
xor2 gate178( .a(N29), .b(N699), .O(N731) );
xor2 gate179( .a(N33), .b(N700), .O(N732) );
xor2 gate180( .a(N37), .b(N701), .O(N733) );
xor2 gate181( .a(N41), .b(N702), .O(N734) );
xor2 gate182( .a(N45), .b(N703), .O(N735) );
xor2 gate183( .a(N49), .b(N704), .O(N736) );
xor2 gate184( .a(N53), .b(N705), .O(N737) );
xor2 gate185( .a(N57), .b(N706), .O(N738) );
xor2 gate186( .a(N61), .b(N707), .O(N739) );
xor2 gate187( .a(N65), .b(N708), .O(N740) );
xor2 gate188( .a(N69), .b(N709), .O(N741) );
xor2 gate189( .a(N73), .b(N710), .O(N742) );
xor2 gate190( .a(N77), .b(N711), .O(N743) );
xor2 gate191( .a(N81), .b(N712), .O(N744) );
xor2 gate192( .a(N85), .b(N713), .O(N745) );
xor2 gate193( .a(N89), .b(N714), .O(N746) );
xor2 gate194( .a(N93), .b(N715), .O(N747) );
xor2 gate195( .a(N97), .b(N716), .O(N748) );
xor2 gate196( .a(N101), .b(N717), .O(N749) );
xor2 gate197( .a(N105), .b(N718), .O(N750) );
xor2 gate198( .a(N109), .b(N719), .O(N751) );
xor2 gate199( .a(N113), .b(N720), .O(N752) );
xor2 gate200( .a(N117), .b(N721), .O(N753) );
xor2 gate201( .a(N121), .b(N722), .O(N754) );
xor2 gate202( .a(N125), .b(N723), .O(N755) );
xor2 gate( .a(X_1), .b(N117_new), .O(N117) );
xor2 gate( .a(X_2), .b(N135_new), .O(N135) );
xor2 gate( .a(X_3), .b(N732), .O(N732_new) );

endmodule