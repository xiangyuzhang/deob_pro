

module c7552 (N1,N5,N9,N12,N15,N18,N23,N26,N29,N32,
              N35,N38,N41,N44,N47,N50,N53,N54,N55,N56,
              N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,
              N69,N70,N73,N74,N75,N76,N77,N78,N79,N80,
              N81,N82,N83,N84,N85,N86,N87,N88,N89,N94,
              N97,N100,N103,N106,N109,N110,N111,N112,N113,N114,
              N115,N118,N121,N124,N127,N130,N133,N134,N135,N138,
              N141,N144,N147,N150,N151,N152,N153,N154,N155,N156,
              N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,
              N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
              N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,
              N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,
              N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
              N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,
              N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,
              N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,
              N237,N238,N239,N240,N242,N245,N248,N251,N254,N257,
              N260,N263,N267,N271,N274,N277,N280,N283,N286,N289,
              N293,N296,N299,N303,N307,N310,N313,N316,N319,N322,
              N325,N328,N331,N334,N337,N340,N343,N346,N349,N352,
              N355,N358,N361,N364,N367,N382,N241_I,N387,N388,N478,
              N482,N484,N486,N489,N492,N501,N505,N507,N509,N511,
              N513,N515,N517,N519,N535,N537,N539,N541,N543,N545,
              N547,N549,N551,N553,N556,N559,N561,N563,N565,N567,
              N569,N571,N573,N582,N643,N707,N813,N881,N882,N883,
              N884,N885,N889,N945,N1110,N1111,N1112,N1113,N1114,N1489,
              N1490,N1781,N10025,N10101,N10102,N10103,N10104,N10109,N10110,N10111,
              N10112,N10350,N10351,N10352,N10353,N10574,N10575,N10576,N10628,N10632,
              N10641,N10704,N10706,N10711,N10712,N10713,N10714,N10715,N10716,N10717,
              N10718,N10729,N10759,N10760,N10761,N10762,N10763,N10827,N10837,N10838,
              N10839,N10840,N10868,N10869,N10870,N10871,N10905,N10906,N10907,N10908,
              N11333,N11334,N11340,N11342,N241_O);

input N1,N5,N9,N12,N15,N18,N23,N26,N29,N32,
      N35,N38,N41,N44,N47,N50,N53,N54,N55,N56,
      N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,
      N69,N70,N73,N74,N75,N76,N77,N78,N79,N80,
      N81,N82,N83,N84,N85,N86,N87,N88,N89,N94,
      N97,N100,N103,N106,N109,N110,N111,N112,N113,N114,
      N115,N118,N121,N124,N127,N130,N133,N134,N135,N138,
      N141,N144,N147,N150,N151,N152,N153,N154,N155,N156,
      N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,
      N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
      N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,
      N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,
      N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
      N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,
      N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,
      N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,
      N237,N238,N239,N240,N242,N245,N248,N251,N254,N257,
      N260,N263,N267,N271,N274,N277,N280,N283,N286,N289,
      N293,N296,N299,N303,N307,N310,N313,N316,N319,N322,
      N325,N328,N331,N334,N337,N340,N343,N346,N349,N352,
      N355,N358,N361,N364,N367,N382,N241_I;

input p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,
        p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,
        p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,
        p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,
        p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,
        p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,
        p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,
        p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,
        p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,
        p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,
        p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,
        p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,
        p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,
        p131,p132,p133,p134,p135,p136,p137,p138,p139,p140,
        p141,p142,p143,p144,p145,p146,p147,p148,p149,p150,
        p151,p152,p153,p154,p155,p156,p157,p158,p159,p160,
        p161,p162,p163,p164,p165,p166,p167,p168,p169,p170,
        p171,p172,p173,p174,p175,p176,p177,p178,p179,p180,
        p181,p182,p183,p184,p185,p186,p187,p188,p189,p190,
        p191,p192,p193,p194,p195,p196,p197,p198,p199,p200,
        p201,p202,p203,p204,p205,p206,p207,p208,p209,p210,
        p211,p212,p213,p214,p215,p216,p217,p218,p219,p220,
        p221,p222,p223,p224,p225,p226,p227,p228,p229,p230,
        p231,p232,p233,p234,p235,p236,p237,p238,p239,p240,
        p241,p242,p243,p244,p245,p246,p247,p248,p249,p250,
        p251,p252,p253,p254,p255,p256,p257,p258,p259,p260,
        p261,p262,p263,p264,p265,p266,p267,p268,p269,p270,
        p271,p272,p273,p274,p275,p276,p277,p278,p279,p280,
        p281,p282,p283,p284,p285,p286,p287,p288,p289,p290,
        p291,p292,p293,p294,p295,p296,p297,p298,p299,p300,
        p301,p302,p303,p304,p305,p306,p307,p308,p309,p310,
        p311,p312,p313,p314,p315,p316,p317,p318,p319,p320,
        p321,p322,p323,p324,p325,p326,p327,p328,p329,p330,
        p331,p332,p333,p334,p335,p336,p337,p338,p339,p340,
        p341,p342,p343,p344,p345,p346,p347,p348,p349,p350,
        p351,p352,p353,p354,p355,p356,p357,p358,p359,p360,
        p361,p362,p363,p364,p365,p366,p367,p368,p369,p370,
        p371,p372,p373,p374,p375,p376,p377,p378,p379,p380,
        p381,p382,p383,p384,p385,p386,p387,p388,p389,p390,
        p391,p392,p393,p394,p395,p396,p397,p398,p399,p400,
        p401,p402,p403,p404,p405,p406,p407,p408,p409,p410,
        p411,p412,p413,p414,p415,p416,p417,p418,p419,p420,
        p421,p422,p423,p424,p425,p426,p427,p428,p429,p430,
        p431,p432,p433,p434,p435,p436,p437,p438,p439,p440,
        p441,p442,p443,p444,p445,p446,p447,p448,p449,p450,
        p451,p452,p453,p454,p455,p456,p457,p458,p459,p460,
        p461,p462,p463,p464,p465,p466,p467,p468,p469,p470,
        p471,p472,p473,p474,p475,p476,p477,p478,p479,p480,
        p481,p482,p483,p484,p485,p486,p487,p488,p489,p490,
        p491,p492,p493,p494,p495,p496,p497,p498,p499,p500,
        p501,p502,p503,p504,p505,p506,p507,p508,p509,p510,
        p511,p512,p513,p514,p515,p516,p517,p518,p519,p520,
        p521,p522,p523,p524,p525,p526,p527,p528,p529,p530,
        p531,p532,p533,p534,p535,p536,p537,p538,p539,p540,
        p541,p542,p543,p544,p545,p546,p547,p548,p549,p550,
        p551,p552,p553,p554,p555,p556,p557,p558,p559,p560,
        p561,p562,p563,p564,p565,p566,p567,p568,p569,p570,
        p571,p572,p573,p574,p575,p576,p577,p578,p579,p580,
        p581,p582,p583,p584,p585,p586,p587,p588,p589,p590,
        p591,p592,p593,p594,p595,p596,p597,p598,p599,p600,
        p601,p602,p603,p604,p605,p606,p607,p608,p609,p610,
        p611,p612,p613,p614,p615,p616,p617,p618,p619,p620,
        p621,p622,p623,p624,p625,p626,p627,p628,p629,p630,
        p631,p632,p633,p634,p635,p636,p637,p638,p639,p640,
        p641,p642,p643,p644,p645,p646,p647,p648,p649,p650,
        p651,p652,p653,p654,p655,p656,p657,p658,p659,p660,
        p661,p662,p663,p664,p665,p666,p667,p668,p669,p670,
        p671,p672,p673,p674,p675,p676,p677,p678,p679,p680,
        p681,p682,p683,p684,p685,p686,p687,p688,p689,p690,
        p691,p692,p693,p694,p695,p696,p697,p698,p699,p700,
        p701,p702,p703,p704,p705,p706,p707,p708,p709,p710,
        p711,p712,p713,p714,p715,p716,p717,p718,p719,p720,
        p721,p722,p723,p724,p725,p726,p727,p728,p729,p730,
        p731,p732,p733,p734,p735,p736,p737,p738,p739,p740,
        p741,p742,p743,p744,p745,p746,p747,p748,p749,p750,
        p751,p752,p753,p754,p755,p756;

output N387,N388,N478,N482,N484,N486,N489,N492,N501,N505,
       N507,N509,N511,N513,N515,N517,N519,N535,N537,N539,
       N541,N543,N545,N547,N549,N551,N553,N556,N559,N561,
       N563,N565,N567,N569,N571,N573,N582,N643,N707,N813,
       N881,N882,N883,N884,N885,N889,N945,N1110,N1111,N1112,
       N1113,N1114,N1489,N1490,N1781,N10025,N10101,N10102,N10103,N10104,
       N10109,N10110,N10111,N10112,N10350,N10351,N10352,N10353,N10574,N10575,
       N10576,N10628,N10632,N10641,N10704,N10706,N10711,N10712,N10713,N10714,
       N10715,N10716,N10717,N10718,N10729,N10759,N10760,N10761,N10762,N10763,
       N10827,N10837,N10838,N10839,N10840,N10868,N10869,N10870,N10871,N10905,
       N10906,N10907,N10908,N11333,N11334,N11340,N11342,N241_O;

wire N467,N469,N494,N528,N575,N578,N585,N590,N593,N596,
     N599,N604,N609,N614,N625,N628,N632,N636,N641,N642,
     N644,N651,N657,N660,N666,N672,N673,N674,N676,N682,
     N688,N689,N695,N700,N705,N706,N708,N715,N721,N727,
     N733,N734,N742,N748,N749,N750,N758,N759,N762,N768,
     N774,N780,N786,N794,N800,N806,N812,N814,N821,N827,
     N833,N839,N845,N853,N859,N865,N871,N886,N887,N957,
     N1028,N1029,N1109,N1115,N1116,N1119,N1125,N1132,N1136,N1141,
     N1147,N1154,N1160,N1167,N1174,N1175,N1182,N1189,N1194,N1199,
     N1206,N1211,N1218,N1222,N1227,N1233,N1240,N1244,N1249,N1256,
     N1263,N1270,N1277,N1284,N1287,N1290,N1293,N1296,N1299,N1302,
     N1305,N1308,N1311,N1314,N1317,N1320,N1323,N1326,N1329,N1332,
     N1335,N1338,N1341,N1344,N1347,N1350,N1353,N1356,N1359,N1362,
     N1365,N1368,N1371,N1374,N1377,N1380,N1383,N1386,N1389,N1392,
     N1395,N1398,N1401,N1404,N1407,N1410,N1413,N1416,N1419,N1422,
     N1425,N1428,N1431,N1434,N1437,N1440,N1443,N1446,N1449,N1452,
     N1455,N1458,N1461,N1464,N1467,N1470,N1473,N1476,N1479,N1482,
     N1485,N1537,N1551,N1649,N1703,N1708,N1713,N1721,N1758,N1782,
     N1783,N1789,N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1805,
     N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,
     N1821,N1822,N1828,N1829,N1830,N1832,N1833,N1834,N1835,N1839,
     N1840,N1841,N1842,N1843,N1845,N1851,N1857,N1858,N1859,N1860,
     N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870,
     N1871,N1872,N1873,N1874,N1875,N1876,N1877,N1878,N1879,N1880,
     N1881,N1882,N1883,N1884,N1885,N1892,N1899,N1906,N1913,N1919,
     N1926,N1927,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,
     N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,N1945,
     N1946,N1947,N1953,N1957,N1958,N1959,N1960,N1961,N1962,N1963,
     N1965,N1966,N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974,
     N1975,N1976,N1977,N1983,N1989,N1990,N1991,N1992,N1993,N1994,
     N1995,N1996,N1997,N2003,N2010,N2011,N2012,N2013,N2014,N2015,
     N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,N2031,
     N2038,N2045,N2052,N2058,N2064,N2065,N2066,N2067,N2068,N2069,
     N2070,N2071,N2072,N2073,N2074,N2081,N2086,N2107,N2108,N2110,
     N2111,N2112,N2113,N2114,N2115,N2117,N2171,N2172,N2230,N2231,
     N2235,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,
     N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,
     N2267,N2268,N2269,N2274,N2275,N2277,N2278,N2279,N2280,N2281,
     N2282,N2283,N2284,N2285,N2286,N2287,N2293,N2299,N2300,N2301,
     N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2315,N2321,
     N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,N2331,
     N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,N2345,N2346,
     N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,
     N2357,N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,
     N2367,N2368,N2374,N2375,N2376,N2377,N2378,N2379,N2380,N2381,
     N2382,N2383,N2384,N2390,N2396,N2397,N2398,N2399,N2400,N2401,
     N2402,N2403,N2404,N2405,N2406,N2412,N2418,N2419,N2420,N2421,
     N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,
     N2432,N2433,N2434,N2435,N2436,N2437,N2441,N2442,N2446,N2450,
     N2454,N2458,N2462,N2466,N2470,N2474,N2478,N2482,N2488,N2496,
     N2502,N2508,N2523,N2533,N2537,N2538,N2542,N2546,N2550,N2554,
     N2561,N2567,N2573,N2604,N2607,N2611,N2615,N2619,N2626,N2632,
     N2638,N2644,N2650,N2653,N2654,N2658,N2662,N2666,N2670,N2674,
     N2680,N2688,N2692,N2696,N2700,N2704,N2728,N2729,N2733,N2737,
     N2741,N2745,N2749,N2753,N2757,N2761,N2765,N2766,N2769,N2772,
     N2775,N2778,N2781,N2784,N2787,N2790,N2793,N2796,N2866,N2867,
     N2868,N2869,N2878,N2913,N2914,N2915,N2916,N2917,N2918,N2919,
     N2920,N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928,N2929,
     N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2988,N3005,
     N3006,N3007,N3008,N3009,N3020,N3021,N3022,N3023,N3024,N3025,
     N3026,N3027,N3028,N3029,N3032,N3033,N3034,N3035,N3036,N3037,
     N3038,N3039,N3040,N3041,N3061,N3064,N3067,N3070,N3073,N3080,
     N3096,N3097,N3101,N3107,N3114,N3122,N3126,N3130,N3131,N3134,
     N3135,N3136,N3137,N3140,N3144,N3149,N3155,N3159,N3167,N3168,
     N3169,N3173,N3178,N3184,N3185,N3189,N3195,N3202,N3210,N3211,
     N3215,N3221,N3228,N3229,N3232,N3236,N3241,N3247,N3251,N3255,
     N3259,N3263,N3267,N3273,N3281,N3287,N3293,N3299,N3303,N3307,
     N3311,N3315,N3322,N3328,N3334,N3340,N3343,N3349,N3355,N3361,
     N3362,N3363,N3364,N3365,N3366,N3367,N3368,N3369,N3370,N3371,
     N3372,N3373,N3374,N3375,N3379,N3380,N3381,N3384,N3390,N3398,
     N3404,N3410,N3416,N3420,N3424,N3428,N3432,N3436,N3440,N3444,
     N3448,N3452,N3453,N3454,N3458,N3462,N3466,N3470,N3474,N3478,
     N3482,N3486,N3487,N3490,N3493,N3496,N3499,N3502,N3507,N3510,
     N3515,N3518,N3521,N3524,N3527,N3530,N3535,N3539,N3542,N3545,
     N3548,N3551,N3552,N3553,N3557,N3560,N3563,N3566,N3569,N3570,
     N3571,N3574,N3577,N3580,N3583,N3586,N3589,N3592,N3595,N3598,
     N3601,N3604,N3607,N3610,N3613,N3616,N3619,N3622,N3625,N3628,
     N3631,N3634,N3637,N3640,N3643,N3646,N3649,N3652,N3655,N3658,
     N3661,N3664,N3667,N3670,N3673,N3676,N3679,N3682,N3685,N3688,
     N3691,N3694,N3697,N3700,N3703,N3706,N3709,N3712,N3715,N3718,
     N3721,N3724,N3727,N3730,N3733,N3736,N3739,N3742,N3745,N3748,
     N3751,N3754,N3757,N3760,N3763,N3766,N3769,N3772,N3775,N3778,
     N3781,N3782,N3783,N3786,N3789,N3792,N3795,N3798,N3801,N3804,
     N3807,N3810,N3813,N3816,N3819,N3822,N3825,N3828,N3831,N3834,
     N3837,N3840,N3843,N3846,N3849,N3852,N3855,N3858,N3861,N3864,
     N3867,N3870,N3873,N3876,N3879,N3882,N3885,N3888,N3891,N3953,
     N3954,N3955,N3956,N3958,N3964,N4193,N4303,N4308,N4313,N4326,
     N4327,N4333,N4334,N4411,N4412,N4463,N4464,N4465,N4466,N4467,
     N4468,N4469,N4470,N4471,N4472,N4473,N4474,N4475,N4476,N4477,
     N4478,N4479,N4480,N4481,N4482,N4483,N4484,N4485,N4486,N4487,
     N4488,N4489,N4490,N4491,N4492,N4493,N4494,N4495,N4496,N4497,
     N4498,N4499,N4500,N4501,N4502,N4503,N4504,N4505,N4506,N4507,
     N4508,N4509,N4510,N4511,N4512,N4513,N4514,N4515,N4516,N4517,
     N4518,N4519,N4520,N4521,N4522,N4523,N4524,N4525,N4526,N4527,
     N4528,N4529,N4530,N4531,N4532,N4533,N4534,N4535,N4536,N4537,
     N4538,N4539,N4540,N4541,N4542,N4543,N4544,N4545,N4549,N4555,
     N4562,N4563,N4566,N4570,N4575,N4576,N4577,N4581,N4586,N4592,
     N4593,N4597,N4603,N4610,N4611,N4612,N4613,N4614,N4615,N4616,
     N4617,N4618,N4619,N4620,N4621,N4622,N4623,N4624,N4625,N4626,
     N4627,N4628,N4629,N4630,N4631,N4632,N4633,N4634,N4635,N4636,
     N4637,N4638,N4639,N4640,N4641,N4642,N4643,N4644,N4645,N4646,
     N4647,N4648,N4649,N4650,N4651,N4652,N4653,N4656,N4657,N4661,
     N4667,N4674,N4675,N4678,N4682,N4687,N4693,N4694,N4695,N4696,
     N4697,N4698,N4699,N4700,N4701,N4702,N4706,N4711,N4717,N4718,
     N4722,N4728,N4735,N4743,N4744,N4745,N4746,N4747,N4748,N4749,
     N4750,N4751,N4752,N4753,N4754,N4755,N4756,N4757,N4758,N4759,
     N4760,N4761,N4762,N4763,N4764,N4765,N4766,N4767,N4768,N4769,
     N4775,N4776,N4777,N4778,N4779,N4780,N4781,N4782,N4783,N4784,
     N4789,N4790,N4793,N4794,N4795,N4796,N4799,N4800,N4801,N4802,
     N4803,N4806,N4809,N4810,N4813,N4814,N4817,N4820,N4823,N4826,
     N4829,N4832,N4835,N4838,N4841,N4844,N4847,N4850,N4853,N4856,
     N4859,N4862,N4865,N4868,N4871,N4874,N4877,N4880,N4883,N4886,
     N4889,N4892,N4895,N4898,N4901,N4904,N4907,N4910,N4913,N4916,
     N4919,N4922,N4925,N4928,N4931,N4934,N4937,N4940,N4943,N4946,
     N4949,N4952,N4955,N4958,N4961,N4964,N4967,N4970,N4973,N4976,
     N4979,N4982,N4985,N4988,N4991,N4994,N4997,N5000,N5003,N5006,
     N5009,N5012,N5015,N5018,N5021,N5024,N5027,N5030,N5033,N5036,
     N5039,N5042,N5045,N5046,N5047,N5048,N5049,N5052,N5055,N5058,
     N5061,N5064,N5065,N5066,N5067,N5068,N5071,N5074,N5077,N5080,
     N5083,N5086,N5089,N5092,N5095,N5098,N5101,N5104,N5107,N5110,
     N5111,N5112,N5113,N5114,N5117,N5120,N5123,N5126,N5129,N5132,
     N5135,N5138,N5141,N5144,N5147,N5150,N5153,N5156,N5159,N5162,
     N5165,N5166,N5167,N5168,N5169,N5170,N5171,N5172,N5173,N5174,
     N5175,N5176,N5177,N5178,N5179,N5180,N5181,N5182,N5183,N5184,
     N5185,N5186,N5187,N5188,N5189,N5190,N5191,N5192,N5193,N5196,
     N5197,N5198,N5199,N5200,N5201,N5202,N5203,N5204,N5205,N5206,
     N5207,N5208,N5209,N5210,N5211,N5212,N5213,N5283,N5284,N5285,
     N5286,N5287,N5288,N5289,N5290,N5291,N5292,N5293,N5294,N5295,
     N5296,N5297,N5298,N5299,N5300,N5314,N5315,N5316,N5317,N5318,
     N5319,N5320,N5321,N5322,N5323,N5324,N5363,N5364,N5365,N5366,
     N5367,N5425,N5426,N5427,N5429,N5430,N5431,N5432,N5433,N5451,
     N5452,N5453,N5454,N5455,N5456,N5457,N5469,N5474,N5475,N5476,
     N5477,N5571,N5572,N5573,N5574,N5584,N5585,N5586,N5587,N5602,
     N5603,N5604,N5605,N5631,N5632,N5640,N5654,N5670,N5683,N5690,
     N5697,N5707,N5718,N5728,N5735,N5736,N5740,N5744,N5747,N5751,
     N5755,N5758,N5762,N5766,N5769,N5770,N5771,N5778,N5789,N5799,
     N5807,N5821,N5837,N5850,N5856,N5863,N5870,N5881,N5892,N5898,
     N5905,N5915,N5926,N5936,N5943,N5944,N5945,N5946,N5947,N5948,
     N5949,N5950,N5951,N5952,N5953,N5954,N5955,N5956,N5957,N5958,
     N5959,N5960,N5966,N5967,N5968,N5969,N5970,N5971,N5972,N5973,
     N5974,N5975,N5976,N5977,N5978,N5979,N5980,N5981,N5989,N5990,
     N5991,N5996,N6000,N6003,N6009,N6014,N6018,N6021,N6022,N6023,
     N6024,N6025,N6026,N6027,N6028,N6029,N6030,N6031,N6032,N6033,
     N6034,N6035,N6036,N6037,N6038,N6039,N6040,N6041,N6047,N6052,
     N6056,N6059,N6060,N6061,N6062,N6063,N6064,N6065,N6066,N6067,
     N6068,N6069,N6070,N6071,N6072,N6073,N6074,N6075,N6076,N6077,
     N6078,N6079,N6083,N6087,N6090,N6091,N6092,N6093,N6094,N6095,
     N6096,N6097,N6098,N6099,N6100,N6101,N6102,N6103,N6104,N6105,
     N6106,N6107,N6108,N6109,N6110,N6111,N6112,N6113,N6114,N6115,
     N6116,N6117,N6118,N6119,N6120,N6121,N6122,N6123,N6124,N6125,
     N6126,N6127,N6131,N6135,N6136,N6137,N6141,N6145,N6148,N6149,
     N6150,N6151,N6152,N6153,N6154,N6155,N6156,N6157,N6158,N6159,
     N6160,N6161,N6162,N6163,N6164,N6165,N6166,N6170,N6174,N6177,
     N6181,N6182,N6183,N6184,N6185,N6186,N6187,N6188,N6189,N6190,
     N6191,N6192,N6193,N6194,N6195,N6196,N6199,N6202,N6203,N6204,
     N6207,N6210,N6213,N6214,N6217,N6220,N6223,N6224,N6225,N6226,
     N6227,N6228,N6229,N6230,N6231,N6232,N6235,N6236,N6239,N6240,
     N6241,N6242,N6243,N6246,N6249,N6252,N6255,N6256,N6257,N6258,
     N6259,N6260,N6261,N6262,N6263,N6266,N6540,N6541,N6542,N6543,
     N6544,N6545,N6546,N6547,N6555,N6556,N6557,N6558,N6559,N6560,
     N6561,N6569,N6594,N6595,N6596,N6597,N6598,N6599,N6600,N6601,
     N6602,N6603,N6604,N6605,N6606,N6621,N6622,N6623,N6624,N6625,
     N6626,N6627,N6628,N6629,N6639,N6640,N6641,N6642,N6643,N6644,
     N6645,N6646,N6647,N6648,N6649,N6650,N6651,N6652,N6653,N6654,
     N6655,N6656,N6657,N6658,N6659,N6660,N6661,N6668,N6677,N6678,
     N6679,N6680,N6681,N6682,N6683,N6684,N6685,N6686,N6687,N6688,
     N6689,N6690,N6702,N6703,N6704,N6705,N6706,N6707,N6708,N6709,
     N6710,N6711,N6712,N6729,N6730,N6731,N6732,N6733,N6734,N6735,
     N6736,N6741,N6742,N6743,N6744,N6751,N6752,N6753,N6754,N6755,
     N6756,N6757,N6758,N6761,N6762,N6766,N6767,N6768,N6769,N6770,
     N6771,N6772,N6773,N6774,N6775,N6776,N6777,N6778,N6779,N6780,
     N6781,N6782,N6783,N6784,N6787,N6788,N6789,N6790,N6791,N6792,
     N6793,N6794,N6795,N6796,N6797,N6800,N6803,N6806,N6809,N6812,
     N6815,N6818,N6821,N6824,N6827,N6830,N6833,N6836,N6837,N6838,
     N6839,N6840,N6841,N6842,N6843,N6844,N6845,N6848,N6849,N6850,
     N6851,N6852,N6853,N6854,N6855,N6856,N6857,N6858,N6859,N6860,
     N6861,N6862,N6863,N6864,N6865,N6866,N6867,N6870,N6871,N6872,
     N6873,N6874,N6875,N6876,N6877,N6878,N6879,N6880,N6881,N6884,
     N6885,N6886,N6887,N6888,N6889,N6890,N6891,N6892,N6893,N6894,
     N6901,N6912,N6923,N6929,N6936,N6946,N6957,N6967,N6968,N6969,
     N6970,N6977,N6988,N6998,N7006,N7020,N7036,N7049,N7055,N7056,
     N7057,N7060,N7061,N7062,N7063,N7064,N7065,N7066,N7067,N7068,
     N7073,N7077,N7080,N7086,N7091,N7095,N7098,N7099,N7100,N7103,
     N7104,N7105,N7106,N7107,N7114,N7125,N7136,N7142,N7149,N7159,
     N7170,N7180,N7187,N7188,N7191,N7194,N7198,N7202,N7205,N7209,
     N7213,N7216,N7219,N7222,N7229,N7240,N7250,N7258,N7272,N7288,
     N7301,N7307,N7314,N7318,N7322,N7325,N7328,N7331,N7334,N7337,
     N7340,N7343,N7346,N7351,N7355,N7358,N7364,N7369,N7373,N7376,
     N7377,N7378,N7381,N7384,N7387,N7391,N7394,N7398,N7402,N7405,
     N7408,N7411,N7414,N7417,N7420,N7423,N7426,N7429,N7432,N7435,
     N7438,N7441,N7444,N7447,N7450,N7453,N7456,N7459,N7462,N7465,
     N7468,N7471,N7474,N7477,N7478,N7479,N7482,N7485,N7488,N7491,
     N7494,N7497,N7500,N7503,N7506,N7509,N7512,N7515,N7518,N7521,
     N7524,N7527,N7530,N7533,N7536,N7539,N7542,N7545,N7548,N7551,
     N7552,N7553,N7556,N7557,N7558,N7559,N7560,N7563,N7566,N7569,
     N7572,N7573,N7574,N7577,N7580,N7581,N7582,N7585,N7588,N7591,
     N7609,N7613,N7620,N7649,N7650,N7655,N7659,N7668,N7671,N7744,
     N7822,N7825,N7826,N7852,N8114,N8117,N8131,N8134,N8144,N8145,
     N8146,N8156,N8166,N8169,N8183,N8186,N8196,N8200,N8204,N8208,
     N8216,N8217,N8218,N8219,N8232,N8233,N8242,N8243,N8244,N8245,
     N8246,N8247,N8248,N8249,N8250,N8251,N8252,N8253,N8254,N8260,
     N8261,N8262,N8269,N8274,N8275,N8276,N8277,N8278,N8279,N8280,
     N8281,N8282,N8283,N8284,N8285,N8288,N8294,N8295,N8296,N8297,
     N8298,N8307,N8315,N8317,N8319,N8321,N8322,N8323,N8324,N8325,
     N8326,N8333,N8337,N8338,N8339,N8340,N8341,N8342,N8343,N8344,
     N8345,N8346,N8347,N8348,N8349,N8350,N8351,N8352,N8353,N8354,
     N8355,N8356,N8357,N8358,N8365,N8369,N8370,N8371,N8372,N8373,
     N8374,N8375,N8376,N8377,N8378,N8379,N8380,N8381,N8382,N8383,
     N8384,N8385,N8386,N8387,N8388,N8389,N8390,N8391,N8392,N8393,
     N8394,N8404,N8405,N8409,N8410,N8411,N8412,N8415,N8416,N8417,
     N8418,N8421,N8430,N8433,N8434,N8435,N8436,N8437,N8438,N8439,
     N8440,N8441,N8442,N8443,N8444,N8447,N8448,N8449,N8450,N8451,
     N8452,N8453,N8454,N8455,N8456,N8457,N8460,N8463,N8466,N8469,
     N8470,N8471,N8474,N8477,N8480,N8483,N8484,N8485,N8488,N8489,
     N8490,N8491,N8492,N8493,N8494,N8495,N8496,N8497,N8500,N8501,
     N8502,N8503,N8504,N8505,N8506,N8507,N8508,N8509,N8510,N8511,
     N8512,N8513,N8514,N8515,N8516,N8517,N8518,N8519,N8522,N8525,
     N8528,N8531,N8534,N8537,N8538,N8539,N8540,N8541,N8545,N8546,
     N8547,N8548,N8551,N8552,N8553,N8554,N8555,N8558,N8561,N8564,
     N8565,N8566,N8569,N8572,N8575,N8578,N8579,N8580,N8583,N8586,
     N8589,N8592,N8595,N8598,N8601,N8604,N8607,N8608,N8609,N8610,
     N8615,N8616,N8617,N8618,N8619,N8624,N8625,N8626,N8627,N8632,
     N8633,N8634,N8637,N8638,N8639,N8644,N8645,N8646,N8647,N8648,
     N8653,N8654,N8655,N8660,N8663,N8666,N8669,N8672,N8675,N8678,
     N8681,N8684,N8687,N8690,N8693,N8696,N8699,N8702,N8705,N8708,
     N8711,N8714,N8717,N8718,N8721,N8724,N8727,N8730,N8733,N8734,
     N8735,N8738,N8741,N8744,N8747,N8750,N8753,N8754,N8755,N8756,
     N8757,N8760,N8763,N8766,N8769,N8772,N8775,N8778,N8781,N8784,
     N8787,N8790,N8793,N8796,N8799,N8802,N8805,N8808,N8811,N8814,
     N8815,N8816,N8817,N8818,N8840,N8857,N8861,N8862,N8863,N8864,
     N8865,N8866,N8871,N8874,N8878,N8879,N8880,N8881,N8882,N8883,
     N8884,N8885,N8886,N8887,N8888,N8898,N8902,N8920,N8924,N8927,
     N8931,N8943,N8950,N8956,N8959,N8960,N8963,N8966,N8991,N8992,
     N8995,N8996,N9001,N9005,N9024,N9025,N9029,N9035,N9053,N9054,
     N9064,N9065,N9066,N9067,N9068,N9071,N9072,N9073,N9074,N9077,
     N9079,N9082,N9083,N9086,N9087,N9088,N9089,N9092,N9093,N9094,
     N9095,N9098,N9099,N9103,N9107,N9111,N9117,N9127,N9146,N9149,
     N9159,N9160,N9161,N9165,N9169,N9173,N9179,N9180,N9181,N9182,
     N9183,N9193,N9203,N9206,N9220,N9223,N9234,N9235,N9236,N9237,
     N9238,N9242,N9243,N9244,N9245,N9246,N9247,N9248,N9249,N9250,
     N9251,N9252,N9256,N9257,N9258,N9259,N9260,N9261,N9262,N9265,
     N9268,N9271,N9272,N9273,N9274,N9275,N9276,N9280,N9285,N9286,
     N9287,N9288,N9290,N9292,N9294,N9296,N9297,N9298,N9299,N9300,
     N9301,N9307,N9314,N9315,N9318,N9319,N9320,N9321,N9322,N9323,
     N9324,N9326,N9332,N9339,N9344,N9352,N9354,N9356,N9358,N9359,
     N9360,N9361,N9362,N9363,N9364,N9365,N9366,N9367,N9368,N9369,
     N9370,N9371,N9372,N9375,N9381,N9382,N9383,N9384,N9385,N9392,
     N9393,N9394,N9395,N9396,N9397,N9398,N9399,N9400,N9401,N9402,
     N9407,N9408,N9412,N9413,N9414,N9415,N9416,N9417,N9418,N9419,
     N9420,N9421,N9422,N9423,N9426,N9429,N9432,N9435,N9442,N9445,
     N9454,N9455,N9456,N9459,N9460,N9461,N9462,N9465,N9466,N9467,
     N9468,N9473,N9476,N9477,N9478,N9485,N9488,N9493,N9494,N9495,
     N9498,N9499,N9500,N9505,N9506,N9507,N9508,N9509,N9514,N9515,
     N9516,N9517,N9520,N9526,N9531,N9539,N9540,N9541,N9543,N9551,
     N9555,N9556,N9557,N9560,N9561,N9562,N9563,N9564,N9565,N9566,
     N9567,N9568,N9569,N9570,N9571,N9575,N9579,N9581,N9582,N9585,
     N9591,N9592,N9593,N9594,N9595,N9596,N9597,N9598,N9599,N9600,
     N9601,N9602,N9603,N9604,N9605,N9608,N9611,N9612,N9613,N9614,
     N9615,N9616,N9617,N9618,N9621,N9622,N9623,N9624,N9626,N9629,
     N9632,N9635,N9642,N9645,N9646,N9649,N9650,N9653,N9656,N9659,
     N9660,N9661,N9662,N9663,N9666,N9667,N9670,N9671,N9674,N9675,
     N9678,N9679,N9682,N9685,N9690,N9691,N9692,N9695,N9698,N9702,
     N9707,N9710,N9711,N9714,N9715,N9716,N9717,N9720,N9721,N9722,
     N9723,N9726,N9727,N9732,N9733,N9734,N9735,N9736,N9737,N9738,
     N9739,N9740,N9741,N9742,N9754,N9758,N9762,N9763,N9764,N9765,
     N9766,N9767,N9768,N9769,N9773,N9774,N9775,N9779,N9784,N9785,
     N9786,N9790,N9791,N9795,N9796,N9797,N9798,N9799,N9800,N9801,
     N9802,N9803,N9805,N9806,N9809,N9813,N9814,N9815,N9816,N9817,
     N9820,N9825,N9826,N9827,N9828,N9829,N9830,N9835,N9836,N9837,
     N9838,N9846,N9847,N9862,N9863,N9866,N9873,N9876,N9890,N9891,
     N9892,N9893,N9894,N9895,N9896,N9897,N9898,N9899,N9900,N9901,
     N9902,N9903,N9904,N9905,N9906,N9907,N9908,N9909,N9910,N9911,
     N9917,N9923,N9924,N9925,N9932,N9935,N9938,N9939,N9945,N9946,
     N9947,N9948,N9949,N9953,N9954,N9955,N9956,N9957,N9958,N9959,
     N9960,N9961,N9964,N9967,N9968,N9969,N9970,N9971,N9972,N9973,
     N9974,N9975,N9976,N9977,N9978,N9979,N9982,N9983,N9986,N9989,
     N9992,N9995,N9996,N9997,N9998,N9999,N10002,N10003,N10006,N10007,
     N10010,N10013,N10014,N10015,N10016,N10017,N10018,N10019,N10020,N10021,
     N10022,N10023,N10024,N10026,N10028,N10032,N10033,N10034,N10035,N10036,
     N10037,N10038,N10039,N10040,N10041,N10042,N10043,N10050,N10053,N10054,
     N10055,N10056,N10057,N10058,N10059,N10060,N10061,N10062,N10067,N10070,
     N10073,N10076,N10077,N10082,N10083,N10084,N10085,N10086,N10093,N10094,
     N10105,N10106,N10107,N10108,N10113,N10114,N10115,N10116,N10119,N10124,
     N10130,N10131,N10132,N10133,N10134,N10135,N10136,N10137,N10138,N10139,
     N10140,N10141,N10148,N10155,N10156,N10157,N10158,N10159,N10160,N10161,
     N10162,N10163,N10164,N10165,N10170,N10173,N10176,N10177,N10178,N10179,
     N10180,N10183,N10186,N10189,N10192,N10195,N10196,N10197,N10200,N10203,
     N10204,N10205,N10206,N10212,N10213,N10230,N10231,N10232,N10233,N10234,
     N10237,N10238,N10239,N10240,N10241,N10242,N10247,N10248,N10259,N10264,
     N10265,N10266,N10267,N10268,N10269,N10270,N10271,N10272,N10273,N10278,
     N10279,N10280,N10281,N10282,N10283,N10287,N10288,N10289,N10290,N10291,
     N10292,N10293,N10294,N10295,N10296,N10299,N10300,N10301,N10306,N10307,
     N10308,N10311,N10314,N10315,N10316,N10317,N10318,N10321,N10324,N10325,
     N10326,N10327,N10328,N10329,N10330,N10331,N10332,N10333,N10334,N10337,
     N10338,N10339,N10340,N10341,N10344,N10354,N10357,N10360,N10367,N10375,
     N10381,N10388,N10391,N10399,N10402,N10406,N10409,N10412,N10415,N10419,
     N10422,N10425,N10428,N10431,N10432,N10437,N10438,N10439,N10440,N10441,
     N10444,N10445,N10450,N10451,N10455,N10456,N10465,N10466,N10479,N10497,
     N10509,N10512,N10515,N10516,N10517,N10518,N10519,N10522,N10525,N10528,
     N10531,N10534,N10535,N10536,N10539,N10542,N10543,N10544,N10545,N10546,
     N10547,N10548,N10549,N10550,N10551,N10552,N10553,N10554,N10555,N10556,
     N10557,N10558,N10559,N10560,N10561,N10562,N10563,N10564,N10565,N10566,
     N10567,N10568,N10569,N10570,N10571,N10572,N10573,N10577,N10581,N10582,
     N10583,N10587,N10588,N10589,N10594,N10595,N10596,N10597,N10598,N10602,
     N10609,N10610,N10621,N10626,N10627,N10629,N10631,N10637,N10638,N10639,
     N10640,N10642,N10643,N10644,N10645,N10647,N10648,N10649,N10652,N10659,
     N10662,N10665,N10668,N10671,N10672,N10673,N10674,N10675,N10678,N10681,
     N10682,N10683,N10684,N10685,N10686,N10687,N10688,N10689,N10690,N10691,
     N10694,N10695,N10696,N10697,N10698,N10701,N10705,N10707,N10708,N10709,
     N10710,N10719,N10720,N10730,N10731,N10737,N10738,N10739,N10746,N10747,
     N10748,N10749,N10750,N10753,N10754,N10764,N10765,N10766,N10767,N10768,
     N10769,N10770,N10771,N10772,N10773,N10774,N10775,N10776,N10778,N10781,
     N10784,N10789,N10792,N10796,N10797,N10798,N10799,N10800,N10803,N10806,
     N10809,N10812,N10815,N10816,N10817,N10820,N10823,N10824,N10825,N10826,
     N10832,N10833,N10834,N10835,N10836,N10845,N10846,N10857,N10862,N10863,
     N10864,N10865,N10866,N10867,N10872,N10873,N10874,N10875,N10876,N10879,
     N10882,N10883,N10884,N10885,N10886,N10887,N10888,N10889,N10890,N10891,
     N10892,N10895,N10896,N10897,N10898,N10899,N10902,N10909,N10910,N10915,
     N10916,N10917,N10918,N10919,N10922,N10923,N10928,N10931,N10934,N10935,
     N10936,N10937,N10938,N10941,N10944,N10947,N10950,N10953,N10954,N10955,
     N10958,N10961,N10962,N10963,N10964,N10969,N10970,N10981,N10986,N10987,
     N10988,N10989,N10990,N10991,N10992,N10995,N10998,N10999,N11000,N11001,
     N11002,N11003,N11004,N11005,N11006,N11007,N11008,N11011,N11012,N11013,
     N11014,N11015,N11018,N11023,N11024,N11027,N11028,N11029,N11030,N11031,
     N11034,N11035,N11040,N11041,N11042,N11043,N11044,N11047,N11050,N11053,
     N11056,N11059,N11062,N11065,N11066,N11067,N11070,N11073,N11074,N11075,
     N11076,N11077,N11078,N11095,N11098,N11099,N11100,N11103,N11106,N11107,
     N11108,N11109,N11110,N11111,N11112,N11113,N11114,N11115,N11116,N11117,
     N11118,N11119,N11120,N11121,N11122,N11123,N11124,N11127,N11130,N11137,
     N11138,N11139,N11140,N11141,N11142,N11143,N11144,N11145,N11152,N11153,
     N11154,N11155,N11156,N11159,N11162,N11165,N11168,N11171,N11174,N11177,
     N11180,N11183,N11184,N11185,N11186,N11187,N11188,N11205,N11210,N11211,
     N11212,N11213,N11214,N11215,N11216,N11217,N11218,N11219,N11220,N11222,
     N11223,N11224,N11225,N11226,N11227,N11228,N11229,N11231,N11232,N11233,
     N11236,N11239,N11242,N11243,N11244,N11245,N11246,N11250,N11252,N11257,
     N11260,N11261,N11262,N11263,N11264,N11265,N11267,N11268,N11269,N11270,
     N11272,N11277,N11278,N11279,N11280,N11282,N11283,N11284,N11285,N11286,
     N11288,N11289,N11290,N11291,N11292,N11293,N11294,N11295,N11296,N11297,
     N11298,N11299,N11302,N11307,N11308,N11309,N11312,N11313,N11314,N11315,
     N11316,N11317,N11320,N11321,N11323,N11327,N11328,N11329,N11331,N11335,
     N11336,N11337,N11338,N11339,N11341,
     N575_NOT,N494_NOT,N957_NOT,N614_NOT,N1029_NOT,N636_NOT,N163_NOT,N1116_NOT,N153_NOT,N1160_NOT,
     N178_NOT,N1175_NOT,N161_NOT,N1182_NOT,N29_NOT,N1211_NOT,N642_NOT,N1249_NOT,N721_NOT,N1270_NOT,
     N727_NOT,N1270_NOT,N734_NOT,N1277_NOT,N1799_NOT,N1814_NOT,N141_NOT,N1845_NOT,N138_NOT,N1845_NOT,
     N135_NOT,N1845_NOT,N141_NOT,N1851_NOT,N135_NOT,N1851_NOT,N124_NOT,N1885_NOT,N103_NOT,N1892_NOT,
     N115_NOT,N1899_NOT,N41_NOT,N1919_NOT,N1947_NOT,N1233_NOT,N77_NOT,N2024_NOT,N79_NOT,N2031_NOT,
     N84_NOT,N2052_NOT,N109_NOT,N2058_NOT,N2239_NOT,N1119_NOT,N2242_NOT,N1119_NOT,N2250_NOT,N1141_NOT,
     N2340_NOT,N1929_NOT,N2349_NOT,N1227_NOT,N2355_NOT,N2172_NOT,N2367_NOT,N1256_NOT,N2436_NOT,N2072_NOT,
     N2354_NOT,N1240_NOT,N2358_NOT,N1989_NOT,N2365_NOT,N1996_NOT,N2257_NOT,N1537_NOT,N202_NOT,N2287_NOT,
     N821_NOT,N2384_NOT,N666_NOT,N2644_NOT,N1167_NOT,N2866_NOT,N660_NOT,N2638_NOT,N651_NOT,N2626_NOT,
     N599_NOT,N2482_NOT,N715_NOT,N2561_NOT,N2918_NOT,N2304_NOT,N2926_NOT,N2324_NOT,N2733_NOT,N2542_NOT,
     N2658_NOT,N2446_NOT,N2488_NOT,N734_NOT,N3070_NOT,N2537_NOT,N2775_NOT,N3569_NOT,N3496_NOT,N1830_NOT,
     N3530_NOT,N1843_NOT,N3652_NOT,N1883_NOT,N806_NOT,N3293_NOT,N859_NOT,N3404_NOT,N3858_NOT,N3486_NOT,
     N4333_NOT,N4334_NOT,N3545_NOT,N4494_NOT,N3563_NOT,N4500_NOT,N1368_NOT,N4536_NOT,N3670_NOT,N4611_NOT,
     N3751_NOT,N4647_NOT,N3754_NOT,N4650_NOT,N3760_NOT,N4652_NOT,N3772_NOT,N4695_NOT,N3798_NOT,N5045_NOT,
     N4481_NOT,N5175_NOT,N5192_NOT,N5193_NOT,N4539_NOT,N5212_NOT,N5316_NOT,N5317_NOT,N5320_NOT,N5321_NOT,
     N4928_NOT,N1973_NOT,N4943_NOT,N4699_NOT,N5049_NOT,N4749_NOT,N1398_NOT,N5957_NOT,N4889_NOT,N6031_NOT,
     N1434_NOT,N6061_NOT,N5117_NOT,N6181_NOT,N5144_NOT,N6187_NOT,N1708_NOT,N6191_NOT,N5640_NOT,N3101_NOT,
     N5654_NOT,N3107_NOT,N5850_NOT,N5789_NOT,N5856_NOT,N5837_NOT,N5870_NOT,N3215_NOT,N3236_NOT,N5915_NOT,
     N6594_NOT,N6024_NOT,N6597_NOT,N6030_NOT,N6105_NOT,N6650_NOT,N6115_NOT,N6655_NOT,N6677_NOT,N6678_NOT,
     N6194_NOT,N6712_NOT,N6743_NOT,N6744_NOT,N3107_NOT,N6782_NOT,N6833_NOT,N6845_NOT,N6977_NOT,N4581_NOT,
     N7057_NOT,N7063_NOT,N3375_NOT,N7100_NOT,N7125_NOT,N4667_NOT,N7258_NOT,N4722_NOT,N7307_NOT,N7288_NOT,
     N3658_NOT,N8323_NOT,N8183_NOT,N6203_NOT,N7574_NOT,N8734_NOT,N7566_NOT,N8756_NOT,N7588_NOT,N8815_NOT,
     N7585_NOT,N8816_NOT,N8864_NOT,N8283_NOT,N7536_NOT,N8881_NOT,N7539_NOT,N8883_NOT,N8672_NOT,N5966_NOT,
     N4193_NOT,N8960_NOT,N8991_NOT,N8483_NOT,N9024_NOT,N8539_NOT,N9053_NOT,N8578_NOT,N9064_NOT,N8608_NOT,
     N9169_NOT,N9356_NOT,N4940_NOT,N9360_NOT,N9368_NOT,N9367_NOT,N9571_NOT,N9301_NOT,N8920_NOT,N9579_NOT,
     N9616_NOT,N9402_NOT,N8950_NOT,N9585_NOT,N8963_NOT,N9591_NOT,N8735_NOT,N9592_NOT,N9029_NOT,N9618_NOT,
     N9623_NOT,N9421_NOT,N5030_NOT,N9715_NOT,N9764_NOT,N9566_NOT,N9765_NOT,N9568_NOT,N9608_NOT,N9375_NOT,
     N8598_NOT,N9899_NOT,N9817_NOT,N9029_NOT,N4871_NOT,N9971_NOT,N9925_NOT,N9895_NOT,N9925_NOT,N9896_NOT,
     N10082_NOT,N9968_NOT,N9478_NOT,N10137_NOT,N7100_NOT,N10140_NOT,N3061_NOT,N10241_NOT,N7620_NOT,N10282_NOT,
     N3241_NOT,N10290_NOT,N9682_NOT,N10332_NOT,N10296_NOT,N4193_NOT,N10439_NOT,N10329_NOT,N10391_NOT,N8950_NOT,
     N5165_NOT,N10367_NOT,N10367_NOT,N3135_NOT,N10381_NOT,N7180_NOT,N9149_NOT,N10534_NOT,N9733_NOT,N10547_NOT,
     N5166_NOT,N10550_NOT,N3159_NOT,N10583_NOT,N10640_NOT,N10564_NOT,N10645_NOT,N10573_NOT,N10709_NOT,N10555_NOT,
     N10652_NOT,N9892_NOT,N10659_NOT,N9245_NOT,N10730_NOT,N10587_NOT,N10753_NOT,N10695_NOT,N7136_NOT,N10784_NOT,
     N10846_NOT,N10799_NOT,N10803_NOT,N8654_NOT,N10820_NOT,N9499_NOT,N8681_NOT,N10886_NOT,N10876_NOT,N8634_NOT,
     N10917_NOT,N10887_NOT,N11029_NOT,N11003_NOT,N7500_NOT,N11042_NOT,N8805_NOT,N11075_NOT,N11056_NOT,N9319_NOT,
     N8778_NOT,N11112_NOT,N7512_NOT,N11118_NOT,N8705_NOT,N11122_NOT,N11130_NOT,N9509_NOT,N8790_NOT,N11185_NOT,
     N7462_NOT,N11215_NOT,N11236_NOT,N9383_NOT,N8796_NOT,N11269_NOT,N11279_NOT,N10283_NOT,N11272_NOT,N9321_NOT,
     N11282_NOT,N11265_NOT,N11312_NOT,N11320_NOT,N11313_NOT,N11321_NOT,N11317_NOT,N11286_NOT,EX1,EX2,EX3,EX4,EX5,EX6,EX7,EX8,EX9,EX10,
     EX11,EX12,EX13,EX14,EX15,EX16,EX17,EX18,EX19,EX20,
     EX21,EX22,EX23,EX24,EX25,EX26,EX27,EX28,EX29,EX30,
     EX31,EX32,EX33,EX34,EX35,EX36,EX37,EX38,EX39,EX40,
     EX41,EX42,EX43,EX44,EX45,EX46,EX47,EX48,EX49,EX50,
     EX51,EX52,EX53,EX54,EX55,EX56,EX57,EX58,EX59,EX60,
     EX61,EX62,EX63,EX64,EX65,EX66,EX67,EX68,EX69,EX70,
     EX71,EX72,EX73,EX74,EX75,EX76,EX77,EX78,EX79,EX80,
     EX81,EX82,EX83,EX84,EX85,EX86,EX87,EX88,EX89,EX90,
     EX91,EX92,EX93,EX94,EX95,EX96,EX97,EX98,EX99,EX100,
     EX101,EX102,EX103,EX104,EX105,EX106,EX107,EX108,EX109,EX110,
     EX111,EX112,EX113,EX114,EX115,EX116,EX117,EX118,EX119,EX120,
     EX121,EX122,EX123,EX124,EX125,EX126,EX127,EX128,EX129,EX130,
     EX131,EX132,EX133,EX134,EX135,EX136,EX137,EX138,EX139,EX140,
     EX141,EX142,EX143,EX144,EX145,EX146,EX147,EX148,EX149,EX150,
     EX151,EX152,EX153,EX154,EX155,EX156,EX157,EX158,EX159,EX160,
     EX161,EX162,EX163,EX164,EX165,EX166,EX167,EX168,EX169,EX170,
     EX171,EX172,EX173,EX174,EX175,EX176,EX177,EX178,EX179,EX180,
     EX181,EX182,EX183,EX184,EX185,EX186,EX187,EX188,EX189,EX190,
     EX191,EX192,EX193,EX194,EX195,EX196,EX197,EX198,EX199,EX200,
     EX201,EX202,EX203,EX204,EX205,EX206,EX207,EX208,EX209,EX210,
     EX211,EX212,EX213,EX214,EX215,EX216,EX217,EX218,EX219,EX220,
     EX221,EX222,EX223,EX224,EX225,EX226,EX227,EX228,EX229,EX230,
     EX231,EX232,EX233,EX234,EX235,EX236,EX237,EX238,EX239,EX240,
     EX241,EX242,EX243,EX244,EX245,EX246,EX247,EX248,EX249,EX250,
     EX251,EX252,EX253,EX254,EX255,EX256,EX257,EX258,EX259,EX260,
     EX261,EX262,EX263,EX264,EX265,EX266,EX267,EX268,EX269,EX270,
     EX271,EX272,EX273,EX274,EX275,EX276,EX277,EX278,EX279,EX280,
     EX281,EX282,EX283,EX284,EX285,EX286,EX287,EX288,EX289,EX290,
     EX291,EX292,EX293,EX294,EX295,EX296,EX297,EX298,EX299,EX300,
     EX301,EX302,EX303,EX304,EX305,EX306,EX307,EX308,EX309,EX310,
     EX311,EX312,EX313,EX314,EX315,EX316,EX317,EX318,EX319,EX320,
     EX321,EX322,EX323,EX324,EX325,EX326,EX327,EX328,EX329,EX330,
     EX331,EX332,EX333,EX334,EX335,EX336,EX337,EX338,EX339,EX340,
     EX341,EX342,EX343,EX344,EX345,EX346,EX347,EX348,EX349,EX350,
     EX351,EX352,EX353,EX354,EX355,EX356,EX357,EX358,EX359,EX360,
     EX361,EX362,EX363,EX364,EX365,EX366,EX367,EX368,EX369,EX370,
     EX371,EX372,EX373,EX374,EX375,EX376,EX377,EX378,EX379,EX380,
     EX381,EX382,EX383,EX384,EX385,EX386,EX387,EX388,EX389,EX390,
     EX391,EX392,EX393,EX394,EX395,EX396,EX397,EX398,EX399,EX400,
     EX401,EX402,EX403,EX404,EX405,EX406,EX407,EX408,EX409,EX410,
     EX411,EX412,EX413,EX414,EX415,EX416,EX417,EX418,EX419,EX420,
     EX421,EX422,EX423,EX424,EX425,EX426,EX427,EX428,EX429,EX430,
     EX431,EX432,EX433,EX434,EX435,EX436,EX437,EX438,EX439,EX440,
     EX441,EX442,EX443,EX444,EX445,EX446,EX447,EX448,EX449,EX450,
     EX451,EX452,EX453,EX454,EX455,EX456,EX457,EX458,EX459,EX460,
     EX461,EX462,EX463,EX464,EX465,EX466,EX467,EX468,EX469,EX470,
     EX471,EX472,EX473,EX474,EX475,EX476,EX477,EX478,EX479,EX480,
     EX481,EX482,EX483,EX484,EX485,EX486,EX487,EX488,EX489,EX490,
     EX491,EX492,EX493,EX494,EX495,EX496,EX497,EX498,EX499,EX500,
     EX501,EX502,EX503,EX504,EX505,EX506,EX507,EX508,EX509,EX510,
     EX511,EX512,EX513,EX514,EX515,EX516,EX517,EX518,EX519,EX520,
     EX521,EX522,EX523,EX524,EX525,EX526,EX527,EX528,EX529,EX530,
     EX531,EX532,EX533,EX534,EX535,EX536,EX537,EX538,EX539,EX540,
     EX541,EX542,EX543,EX544,EX545,EX546,EX547,EX548,EX549,EX550,
     EX551,EX552,EX553,EX554,EX555,EX556,EX557,EX558,EX559,EX560,
     EX561,EX562,EX563,EX564,EX565,EX566,EX567,EX568,EX569,EX570,
     EX571,EX572,EX573,EX574,EX575,EX576,EX577,EX578,EX579,EX580,
     EX581,EX582,EX583,EX584,EX585,EX586,EX587,EX588,EX589,EX590,
     EX591,EX592,EX593,EX594,EX595,EX596,EX597,EX598,EX599,EX600,
     EX601,EX602,EX603,EX604,EX605,EX606,EX607,EX608,EX609,EX610,
     EX611,EX612,EX613,EX614,EX615,EX616,EX617,EX618,EX619,EX620,
     EX621,EX622,EX623,EX624,EX625,EX626,EX627,EX628,EX629,EX630,
     EX631,EX632,EX633,EX634,EX635,EX636,EX637,EX638,EX639,EX640,
     EX641,EX642,EX643,EX644,EX645,EX646,EX647,EX648,EX649,EX650,
     EX651,EX652,EX653,EX654,EX655,EX656,EX657,EX658,EX659,EX660,
     EX661,EX662,EX663,EX664,EX665,EX666,EX667,EX668,EX669,EX670,
     EX671,EX672,EX673,EX674,EX675,EX676,EX677,EX678,EX679,EX680,
     EX681,EX682,EX683,EX684,EX685,EX686,EX687,EX688,EX689,EX690,
     EX691,EX692,EX693,EX694,EX695,EX696,EX697,EX698,EX699,EX700,
     EX701,EX702,EX703,EX704,EX705,EX706,EX707,EX708,EX709,EX710,
     EX711,EX712,EX713,EX714,EX715,EX716,EX717,EX718,EX719,EX720,
     EX721,EX722,EX723,EX724,EX725,EX726,EX727,EX728,EX729,EX730,
     EX731,EX732,EX733,EX734,EX735,EX736,EX737,EX738,EX739,EX740,
     EX741,EX742,EX743,EX744,EX745,EX746,EX747,EX748,EX749,EX750,
     EX751,EX752,EX753,EX754,EX755,EX756,EX757,EX758,EX759,EX760,
     EX761,EX762,EX763,EX764,EX765,EX766,EX767,EX768,EX769,EX770,
     EX771,EX772,EX773,EX774,EX775,EX776,EX777,EX778,EX779,EX780,
     EX781,EX782,EX783,EX784,EX785,EX786,EX787,EX788,EX789,EX790,
     EX791,EX792,EX793,EX794,EX795,EX796,EX797,EX798,EX799,EX800,
     EX801,EX802,EX803,EX804,EX805,EX806,EX807,EX808,EX809,EX810,
     EX811,EX812,EX813,EX814,EX815,EX816,EX817,EX818,EX819,EX820,
     EX821,EX822,EX823,EX824,EX825,EX826,EX827,EX828,EX829,EX830,
     EX831,EX832,EX833,EX834,EX835,EX836,EX837,EX838,EX839,EX840,
     EX841,EX842,EX843,EX844,EX845,EX846,EX847,EX848,EX849,EX850,
     EX851,EX852,EX853,EX854,EX855,EX856,EX857,EX858,EX859,EX860,
     EX861,EX862,EX863,EX864,EX865,EX866,EX867,EX868,EX869,EX870,
     EX871,EX872,EX873,EX874,EX875,EX876,EX877,EX878,EX879,EX880,
     EX881,EX882,EX883,EX884,EX885,EX886,EX887,EX888,EX889,EX890,
     EX891,EX892,EX893,EX894,EX895,EX896,EX897,EX898,EX899,EX900,
     EX901,EX902,EX903,EX904,EX905,EX906,EX907,EX908,EX909,EX910,
     EX911,EX912,EX913,EX914,EX915,EX916,EX917,EX918,EX919,EX920,
     EX921,EX922,EX923,EX924,EX925,EX926,EX927,EX928,EX929,EX930,
     EX931,EX932,EX933,EX934,EX935,EX936,EX937,EX938,EX939,EX940,
     EX941,EX942,EX943,EX944,EX945,EX946,EX947,EX948,EX949,EX950,
     EX951,EX952,EX953,EX954,EX955,EX956,EX957,EX958,EX959,EX960,
     EX961,EX962,EX963,EX964,EX965,EX966,EX967,EX968,EX969,EX970,
     EX971,EX972,EX973,EX974,EX975,EX976,EX977,EX978,EX979,EX980,
     EX981,EX982,EX983,EX984,EX985,EX986,EX987,EX988,EX989,EX990,
     EX991,EX992,EX993,EX994,EX995,EX996,EX997,EX998,EX999,EX1000,
     EX1001,EX1002,EX1003,EX1004,EX1005,EX1006,EX1007,EX1008,EX1009,EX1010,
     EX1011,EX1012,EX1013,EX1014,EX1015,EX1016,EX1017,EX1018,EX1019,EX1020,
     EX1021,EX1022,EX1023,EX1024,EX1025,EX1026,EX1027,EX1028,EX1029,EX1030,
     EX1031,EX1032,EX1033,EX1034,EX1035,EX1036,EX1037,EX1038,EX1039,EX1040,
     EX1041,EX1042,EX1043,EX1044,EX1045,EX1046,EX1047,EX1048,EX1049,EX1050,
     EX1051,EX1052,EX1053,EX1054,EX1055,EX1056,EX1057,EX1058,EX1059,EX1060,
     EX1061,EX1062,EX1063,EX1064,EX1065,EX1066,EX1067,EX1068,EX1069,EX1070,
     EX1071,EX1072,EX1073,EX1074,EX1075,EX1076,EX1077,EX1078,EX1079,EX1080,
     EX1081,EX1082,EX1083,EX1084,EX1085,EX1086,EX1087,EX1088,EX1089,EX1090,
     EX1091,EX1092,EX1093,EX1094,EX1095,EX1096,EX1097,EX1098,EX1099,EX1100,
     EX1101,EX1102,EX1103,EX1104,EX1105,EX1106,EX1107,EX1108,EX1109,EX1110,
     EX1111,EX1112,EX1113,EX1114,EX1115,EX1116,EX1117,EX1118,EX1119,EX1120,
     EX1121,EX1122,EX1123,EX1124,EX1125,EX1126,EX1127,EX1128,EX1129,EX1130,
     EX1131,EX1132,EX1133,EX1134,EX1135,EX1136,EX1137,EX1138,EX1139,EX1140,
     EX1141,EX1142,EX1143,EX1144,EX1145,EX1146,EX1147,EX1148,EX1149,EX1150,
     EX1151,EX1152,EX1153,EX1154,EX1155,EX1156,EX1157,EX1158,EX1159,EX1160,
     EX1161,EX1162,EX1163,EX1164,EX1165,EX1166,EX1167,EX1168,EX1169,EX1170,
     EX1171,EX1172,EX1173,EX1174,EX1175,EX1176,EX1177,EX1178,EX1179,EX1180,
     EX1181,EX1182,EX1183,EX1184,EX1185,EX1186,EX1187,EX1188,EX1189,EX1190,
     EX1191,EX1192,EX1193,EX1194,EX1195,EX1196,EX1197,EX1198,EX1199,EX1200,
     EX1201,EX1202,EX1203,EX1204,EX1205,EX1206,EX1207,EX1208,EX1209,EX1210,
     EX1211,EX1212,EX1213,EX1214,EX1215,EX1216,EX1217,EX1218,EX1219,EX1220,
     EX1221,EX1222,EX1223,EX1224,EX1225,EX1226,EX1227,EX1228,EX1229,EX1230,
     EX1231,EX1232,EX1233,EX1234,EX1235,EX1236,EX1237,EX1238,EX1239,EX1240,
     EX1241,EX1242,EX1243,EX1244,EX1245,EX1246,EX1247,EX1248,EX1249,EX1250,
     EX1251,EX1252,EX1253,EX1254,EX1255,EX1256,EX1257,EX1258,EX1259,EX1260,
     EX1261,EX1262,EX1263,EX1264,EX1265,EX1266,EX1267,EX1268,EX1269,EX1270,
     EX1271,EX1272,EX1273,EX1274,EX1275,EX1276,EX1277,EX1278,EX1279,EX1280,
     EX1281,EX1282,EX1283,EX1284,EX1285,EX1286,EX1287,EX1288,EX1289,EX1290,
     EX1291,EX1292,EX1293,EX1294,EX1295,EX1296,EX1297,EX1298,EX1299,EX1300,
     EX1301,EX1302,EX1303,EX1304,EX1305,EX1306,EX1307,EX1308,EX1309,EX1310,
     EX1311,EX1312,EX1313,EX1314,EX1315,EX1316,EX1317,EX1318,EX1319,EX1320,
     EX1321,EX1322,EX1323,EX1324,EX1325,EX1326,EX1327,EX1328,EX1329,EX1330,
     EX1331,EX1332,EX1333,EX1334,EX1335,EX1336,EX1337,EX1338,EX1339,EX1340,
     EX1341,EX1342,EX1343,EX1344,EX1345,EX1346,EX1347,EX1348,EX1349,EX1350,
     EX1351,EX1352,EX1353,EX1354,EX1355,EX1356,EX1357,EX1358,EX1359,EX1360,
     EX1361,EX1362,EX1363,EX1364,EX1365,EX1366,EX1367,EX1368,EX1369,EX1370,
     EX1371,EX1372,EX1373,EX1374,EX1375,EX1376,EX1377,EX1378,EX1379,EX1380,
     EX1381,EX1382,EX1383,EX1384,EX1385,EX1386,EX1387,EX1388,EX1389,EX1390,
     EX1391,EX1392,EX1393,EX1394,EX1395,EX1396,EX1397,EX1398,EX1399,EX1400,
     EX1401,EX1402,EX1403,EX1404,EX1405,EX1406,EX1407,EX1408,EX1409,EX1410,
     EX1411,EX1412,EX1413,EX1414,EX1415,EX1416,EX1417,EX1418,EX1419,EX1420,
     EX1421,EX1422,EX1423,EX1424,EX1425,EX1426,EX1427,EX1428,EX1429,EX1430,
     EX1431,EX1432,EX1433,EX1434,EX1435,EX1436,EX1437,EX1438,EX1439,EX1440,
     EX1441,EX1442,EX1443,EX1444,EX1445,EX1446,EX1447,EX1448,EX1449,EX1450,
     EX1451,EX1452,EX1453,EX1454,EX1455,EX1456,EX1457,EX1458,EX1459,EX1460,
     EX1461,EX1462,EX1463,EX1464,EX1465,EX1466,EX1467,EX1468,EX1469,EX1470,
     EX1471,EX1472,EX1473,EX1474,EX1475,EX1476,EX1477,EX1478,EX1479,EX1480,
     EX1481,EX1482,EX1483,EX1484,EX1485,EX1486,EX1487,EX1488,EX1489,EX1490,
     EX1491,EX1492,EX1493,EX1494,EX1495,EX1496,EX1497,EX1498,EX1499,EX1500,
     EX1501,EX1502,EX1503,EX1504,EX1505,EX1506,EX1507,EX1508,EX1509,EX1510,
     EX1511,EX1512,EX1513,EX1514,EX1515,EX1516,EX1517,EX1518,EX1519,EX1520,
     EX1521,EX1522,EX1523,EX1524,EX1525,EX1526,EX1527,EX1528,EX1529,EX1530,
     EX1531,EX1532,EX1533,EX1534,EX1535,EX1536,EX1537,EX1538,EX1539,EX1540,
     EX1541,EX1542,EX1543,EX1544,EX1545,EX1546,EX1547,EX1548,EX1549,EX1550,
     EX1551,EX1552,EX1553,EX1554,EX1555,EX1556,EX1557,EX1558,EX1559,EX1560,
     EX1561,EX1562,EX1563,EX1564,EX1565,EX1566,EX1567,EX1568,EX1569,EX1570,
     EX1571,EX1572,EX1573,EX1574,EX1575,EX1576,EX1577,EX1578,EX1579,EX1580,
     EX1581,EX1582,EX1583,EX1584,EX1585,EX1586,EX1587,EX1588,EX1589,EX1590,
     EX1591,EX1592,EX1593,EX1594,EX1595,EX1596,EX1597,EX1598,EX1599,EX1600,
     EX1601,EX1602,EX1603,EX1604,EX1605,EX1606,EX1607,EX1608,EX1609,EX1610,
     EX1611,EX1612,EX1613,EX1614,EX1615,EX1616,EX1617,EX1618,EX1619,EX1620,
     EX1621,EX1622,EX1623,EX1624,EX1625,EX1626,EX1627,EX1628,EX1629,EX1630,
     EX1631,EX1632,EX1633,EX1634,EX1635,EX1636,EX1637,EX1638,EX1639,EX1640,
     EX1641,EX1642,EX1643,EX1644,EX1645,EX1646,EX1647,EX1648,EX1649,EX1650,
     EX1651,EX1652,EX1653,EX1654,EX1655,EX1656,EX1657,EX1658,EX1659,EX1660,
     EX1661,EX1662,EX1663,EX1664,EX1665,EX1666,EX1667,EX1668,EX1669,EX1670,
     EX1671,EX1672,EX1673,EX1674,EX1675,EX1676,EX1677,EX1678,EX1679,EX1680,
     EX1681,EX1682,EX1683,EX1684,EX1685,EX1686,EX1687,EX1688,EX1689,EX1690,
     EX1691,EX1692,EX1693,EX1694,EX1695,EX1696,EX1697,EX1698,EX1699,EX1700,
     EX1701,EX1702,EX1703,EX1704,EX1705,EX1706,EX1707,EX1708,EX1709,EX1710,
     EX1711,EX1712,EX1713,EX1714,EX1715,EX1716,EX1717,EX1718,EX1719,EX1720,
     EX1721,EX1722,EX1723,EX1724,EX1725,EX1726,EX1727,EX1728,EX1729,EX1730,
     EX1731,EX1732,EX1733,EX1734,EX1735,EX1736,EX1737,EX1738,EX1739,EX1740,
     EX1741,EX1742,EX1743,EX1744,EX1745,EX1746,EX1747,EX1748,EX1749,EX1750,
     EX1751,EX1752,EX1753,EX1754,EX1755,EX1756,EX1757,EX1758,EX1759,EX1760,
     EX1761,EX1762,EX1763,EX1764,EX1765,EX1766,EX1767,EX1768,EX1769,EX1770,
     EX1771,EX1772,EX1773,EX1774,EX1775,EX1776,EX1777,EX1778,EX1779,EX1780,
     EX1781,EX1782,EX1783,EX1784,EX1785,EX1786,EX1787,EX1788,EX1789,EX1790,
     EX1791,EX1792,EX1793,EX1794,EX1795,EX1796,EX1797,EX1798,EX1799,EX1800,
     EX1801,EX1802,EX1803,EX1804,EX1805,EX1806,EX1807,EX1808,EX1809,EX1810,
     EX1811,EX1812,EX1813,EX1814,EX1815,EX1816,EX1817,EX1818,EX1819,EX1820,
     EX1821,EX1822,EX1823,EX1824,EX1825,EX1826,EX1827,EX1828,EX1829,EX1830,
     EX1831,EX1832,EX1833,EX1834,EX1835,EX1836,EX1837,EX1838,EX1839,EX1840,
     EX1841,EX1842,EX1843,EX1844,EX1845,EX1846,EX1847,EX1848,EX1849,EX1850,
     EX1851,EX1852,EX1853,EX1854,EX1855,EX1856,EX1857,EX1858,EX1859,EX1860,
     EX1861,EX1862,EX1863,EX1864,EX1865,EX1866,EX1867,EX1868,EX1869,EX1870,
     EX1871,EX1872,EX1873,EX1874,EX1875,EX1876,EX1877,EX1878,EX1879,EX1880,
     EX1881,EX1882,EX1883,EX1884,EX1885,EX1886,EX1887,EX1888,EX1889,EX1890;


buf1 gate1( .a(N1), .O(N387) );
buf1 gate2( .a(N1), .O(N388) );
inv1 gate3( .a(N57), .O(N467) );
and2 gate4( .a(N134), .b(N133), .O(N469) );
buf1 gate5( .a(N248), .O(N478) );
buf1 gate6( .a(N254), .O(N482) );
buf1 gate7( .a(N257), .O(N484) );
buf1 gate8( .a(N260), .O(N486) );
buf1 gate9( .a(N263), .O(N489) );
buf1 gate10( .a(N267), .O(N492) );
and4 gate11( .a(N162), .b(N172), .c(N188), .d(N199), .O(N494) );
buf1 gate12( .a(N274), .O(N501) );
buf1 gate13( .a(N280), .O(N505) );
buf1 gate14( .a(N283), .O(N507) );
buf1 gate15( .a(N286), .O(N509) );
buf1 gate16( .a(N289), .O(N511) );
buf1 gate17( .a(N293), .O(N513) );
buf1 gate18( .a(N296), .O(N515) );
buf1 gate19( .a(N299), .O(N517) );
buf1 gate20( .a(N303), .O(N519) );
and4 gate21( .a(N150), .b(N184), .c(N228), .d(N240), .O(N528) );
buf1 gate22( .a(N307), .O(N535) );
buf1 gate23( .a(N310), .O(N537) );
buf1 gate24( .a(N313), .O(N539) );
buf1 gate25( .a(N316), .O(N541) );
buf1 gate26( .a(N319), .O(N543) );
buf1 gate27( .a(N322), .O(N545) );
buf1 gate28( .a(N325), .O(N547) );
buf1 gate29( .a(N328), .O(N549) );
buf1 gate30( .a(N331), .O(N551) );
buf1 gate31( .a(N334), .O(N553) );
buf1 gate32( .a(N337), .O(N556) );
buf1 gate33( .a(N343), .O(N559) );
buf1 gate34( .a(N346), .O(N561) );
buf1 gate35( .a(N349), .O(N563) );
buf1 gate36( .a(N352), .O(N565) );
buf1 gate37( .a(N355), .O(N567) );
buf1 gate38( .a(N358), .O(N569) );
buf1 gate39( .a(N361), .O(N571) );
buf1 gate40( .a(N364), .O(N573) );
and4 gate41( .a(N183), .b(N182), .c(N185), .d(N186), .O(N575) );
and4 gate42( .a(N210), .b(N152), .c(N218), .d(N230), .O(N578) );
inv1 gate43( .a(N15), .O(N582) );
inv1 gate44( .a(N5), .O(N585) );
buf1 gate45( .a(N1), .O(N590) );
inv1 gate46( .a(N5), .O(N593) );
inv1 gate47( .a(N5), .O(N596) );
inv1 gate48( .a(N289), .O(N599) );
inv1 gate49( .a(N299), .O(N604) );
inv1 gate50( .a(N303), .O(N609) );
buf1 gate51( .a(N38), .O(N614) );
buf1 gate52( .a(N15), .O(N625) );
nand2 gate53( .a(N12), .b(N9), .O(N628) );
nand2 gate54( .a(N12), .b(N9), .O(N632) );
buf1 gate55( .a(N38), .O(N636) );
inv1 gate56( .a(N245), .O(N641) );
inv1 gate57( .a(N248), .O(N642) );
buf1 gate58( .a(N251), .O(N643) );
inv1 gate59( .a(N251), .O(N644) );
inv1 gate60( .a(N254), .O(N651) );
buf1 gate61( .a(N106), .O(N657) );
inv1 gate62( .a(N257), .O(N660) );
inv1 gate63( .a(N260), .O(N666) );
inv1 gate64( .a(N263), .O(N672) );
inv1 gate65( .a(N267), .O(N673) );
inv1 gate66( .a(N106), .O(N674) );
buf1 gate67( .a(N18), .O(N676) );
buf1 gate68( .a(N18), .O(N682) );
and2 gate69( .a(N382), .b(N263), .O(N688) );
buf1 gate70( .a(N18), .O(N689) );
inv1 gate71( .a(N18), .O(N695) );
nand2 gate72( .a(N382), .b(N267), .O(N700) );
inv1 gate73( .a(N271), .O(N705) );
inv1 gate74( .a(N274), .O(N706) );
buf1 gate75( .a(N277), .O(N707) );
inv1 gate76( .a(N277), .O(N708) );
inv1 gate77( .a(N280), .O(N715) );
inv1 gate78( .a(N283), .O(N721) );
inv1 gate79( .a(N286), .O(N727) );
inv1 gate80( .a(N289), .O(N733) );
inv1 gate81( .a(N293), .O(N734) );
inv1 gate82( .a(N296), .O(N742) );
inv1 gate83( .a(N299), .O(N748) );
inv1 gate84( .a(N303), .O(N749) );
buf1 gate85( .a(N367), .O(N750) );
inv1 gate86( .a(N307), .O(N758) );
inv1 gate87( .a(N310), .O(N759) );
inv1 gate88( .a(N313), .O(N762) );
inv1 gate89( .a(N316), .O(N768) );
inv1 gate90( .a(N319), .O(N774) );
inv1 gate91( .a(N322), .O(N780) );
inv1 gate92( .a(N325), .O(N786) );
inv1 gate93( .a(N328), .O(N794) );
inv1 gate94( .a(N331), .O(N800) );
inv1 gate95( .a(N334), .O(N806) );
inv1 gate96( .a(N337), .O(N812) );
buf1 gate97( .a(N340), .O(N813) );
inv1 gate98( .a(N340), .O(N814) );
inv1 gate99( .a(N343), .O(N821) );
inv1 gate100( .a(N346), .O(N827) );
inv1 gate101( .a(N349), .O(N833) );
inv1 gate102( .a(N352), .O(N839) );
inv1 gate103( .a(N355), .O(N845) );
inv1 gate104( .a(N358), .O(N853) );
inv1 gate105( .a(N361), .O(N859) );
inv1 gate106( .a(N364), .O(N865) );
buf1 gate107( .a(N367), .O(N871) );
nand2 gate108( .a(N467), .b(N585), .O(N881) );
inv1 gate109( .a(N528), .O(N882) );
inv1 gate110( .a(N578), .O(N883) );
inv1 gate111( .a(N575), .O(N884) );
inv1 gate112( .a(N494), .O(N885) );
and2 gate113( .a(N528), .b(N578), .O(N886) );
inv1 gate( .a(N575),.O(N575_NOT) );
inv1 gate( .a(N494),.O(N494_NOT));
and2 gate( .a(N575_NOT), .b(p1), .O(EX1) );
and2 gate( .a(N494_NOT), .b(EX1), .O(EX2) );
and2 gate( .a(N575), .b(p2), .O(EX3) );
and2 gate( .a(N494_NOT), .b(EX3), .O(EX4) );
and2 gate( .a(N575_NOT), .b(p3), .O(EX5) );
and2 gate( .a(N494), .b(EX5), .O(EX6) );
and2 gate( .a(N575), .b(p4), .O(EX7) );
and2 gate( .a(N494), .b(EX7), .O(EX8) );
or2  gate( .a(EX2), .b(EX4), .O(EX9) );
or2  gate( .a(EX6), .b(EX9), .O(EX10) );
or2  gate( .a(EX8), .b(EX10), .O(N887) );
buf1 gate115( .a(N590), .O(N889) );
buf1 gate116( .a(N657), .O(N945) );
inv1 gate117( .a(N688), .O(N957) );
and2 gate118( .a(N382), .b(N641), .O(N1028) );
nand2 gate119( .a(N382), .b(N705), .O(N1029) );
and2 gate120( .a(N469), .b(N596), .O(N1109) );
nand2 gate121( .a(N242), .b(N593), .O(N1110) );
inv1 gate122( .a(N625), .O(N1111) );
nand2 gate123( .a(N242), .b(N593), .O(N1112) );
nand2 gate124( .a(N469), .b(N596), .O(N1113) );
inv1 gate125( .a(N625), .O(N1114) );
inv1 gate126( .a(N871), .O(N1115) );
buf1 gate127( .a(N590), .O(N1116) );
buf1 gate128( .a(N628), .O(N1119) );
buf1 gate129( .a(N682), .O(N1125) );
buf1 gate130( .a(N628), .O(N1132) );
buf1 gate131( .a(N682), .O(N1136) );
buf1 gate132( .a(N628), .O(N1141) );
buf1 gate133( .a(N682), .O(N1147) );
buf1 gate134( .a(N632), .O(N1154) );
buf1 gate135( .a(N676), .O(N1160) );
and2 gate136( .a(N700), .b(N614), .O(N1167) );
and2 gate137( .a(N700), .b(N614), .O(N1174) );
buf1 gate138( .a(N682), .O(N1175) );
buf1 gate139( .a(N676), .O(N1182) );
inv1 gate140( .a(N657), .O(N1189) );
inv1 gate141( .a(N676), .O(N1194) );
inv1 gate142( .a(N682), .O(N1199) );
inv1 gate143( .a(N689), .O(N1206) );
buf1 gate144( .a(N695), .O(N1211) );
inv1 gate145( .a(N750), .O(N1218) );
inv1 gate146( .a(N1028), .O(N1222) );
buf1 gate147( .a(N632), .O(N1227) );
buf1 gate148( .a(N676), .O(N1233) );
buf1 gate149( .a(N632), .O(N1240) );
buf1 gate150( .a(N676), .O(N1244) );
buf1 gate151( .a(N689), .O(N1249) );
buf1 gate152( .a(N689), .O(N1256) );
buf1 gate153( .a(N695), .O(N1263) );
buf1 gate154( .a(N689), .O(N1270) );
buf1 gate155( .a(N689), .O(N1277) );
buf1 gate156( .a(N700), .O(N1284) );
buf1 gate157( .a(N614), .O(N1287) );
buf1 gate158( .a(N666), .O(N1290) );
buf1 gate159( .a(N660), .O(N1293) );
buf1 gate160( .a(N651), .O(N1296) );
buf1 gate161( .a(N614), .O(N1299) );
buf1 gate162( .a(N644), .O(N1302) );
buf1 gate163( .a(N700), .O(N1305) );
buf1 gate164( .a(N614), .O(N1308) );
buf1 gate165( .a(N614), .O(N1311) );
buf1 gate166( .a(N666), .O(N1314) );
buf1 gate167( .a(N660), .O(N1317) );
buf1 gate168( .a(N651), .O(N1320) );
buf1 gate169( .a(N644), .O(N1323) );
buf1 gate170( .a(N609), .O(N1326) );
buf1 gate171( .a(N604), .O(N1329) );
buf1 gate172( .a(N742), .O(N1332) );
buf1 gate173( .a(N599), .O(N1335) );
buf1 gate174( .a(N727), .O(N1338) );
buf1 gate175( .a(N721), .O(N1341) );
buf1 gate176( .a(N715), .O(N1344) );
buf1 gate177( .a(N734), .O(N1347) );
buf1 gate178( .a(N708), .O(N1350) );
buf1 gate179( .a(N609), .O(N1353) );
buf1 gate180( .a(N604), .O(N1356) );
buf1 gate181( .a(N742), .O(N1359) );
buf1 gate182( .a(N734), .O(N1362) );
buf1 gate183( .a(N599), .O(N1365) );
buf1 gate184( .a(N727), .O(N1368) );
buf1 gate185( .a(N721), .O(N1371) );
buf1 gate186( .a(N715), .O(N1374) );
buf1 gate187( .a(N708), .O(N1377) );
buf1 gate188( .a(N806), .O(N1380) );
buf1 gate189( .a(N800), .O(N1383) );
buf1 gate190( .a(N794), .O(N1386) );
buf1 gate191( .a(N786), .O(N1389) );
buf1 gate192( .a(N780), .O(N1392) );
buf1 gate193( .a(N774), .O(N1395) );
buf1 gate194( .a(N768), .O(N1398) );
buf1 gate195( .a(N762), .O(N1401) );
buf1 gate196( .a(N806), .O(N1404) );
buf1 gate197( .a(N800), .O(N1407) );
buf1 gate198( .a(N794), .O(N1410) );
buf1 gate199( .a(N780), .O(N1413) );
buf1 gate200( .a(N774), .O(N1416) );
buf1 gate201( .a(N768), .O(N1419) );
buf1 gate202( .a(N762), .O(N1422) );
buf1 gate203( .a(N786), .O(N1425) );
buf1 gate204( .a(N636), .O(N1428) );
buf1 gate205( .a(N636), .O(N1431) );
buf1 gate206( .a(N865), .O(N1434) );
buf1 gate207( .a(N859), .O(N1437) );
buf1 gate208( .a(N853), .O(N1440) );
buf1 gate209( .a(N845), .O(N1443) );
buf1 gate210( .a(N839), .O(N1446) );
buf1 gate211( .a(N833), .O(N1449) );
buf1 gate212( .a(N827), .O(N1452) );
buf1 gate213( .a(N821), .O(N1455) );
buf1 gate214( .a(N814), .O(N1458) );
buf1 gate215( .a(N865), .O(N1461) );
buf1 gate216( .a(N859), .O(N1464) );
buf1 gate217( .a(N853), .O(N1467) );
buf1 gate218( .a(N839), .O(N1470) );
buf1 gate219( .a(N833), .O(N1473) );
buf1 gate220( .a(N827), .O(N1476) );
buf1 gate221( .a(N821), .O(N1479) );
buf1 gate222( .a(N845), .O(N1482) );
buf1 gate223( .a(N814), .O(N1485) );
inv1 gate224( .a(N1109), .O(N1489) );
buf1 gate225( .a(N1116), .O(N1490) );
inv1 gate( .a(N957),.O(N957_NOT) );
inv1 gate( .a(N614),.O(N614_NOT));
and2 gate( .a(N957_NOT), .b(p5), .O(EX11) );
and2 gate( .a(N614_NOT), .b(EX11), .O(EX12) );
and2 gate( .a(N957), .b(p6), .O(EX13) );
and2 gate( .a(N614_NOT), .b(EX13), .O(EX14) );
and2 gate( .a(N957_NOT), .b(p7), .O(EX15) );
and2 gate( .a(N614), .b(EX15), .O(EX16) );
and2 gate( .a(N957), .b(p8), .O(EX17) );
and2 gate( .a(N614), .b(EX17), .O(EX18) );
or2  gate( .a(EX12), .b(EX14), .O(EX19) );
or2  gate( .a(EX16), .b(EX19), .O(EX20) );
or2  gate( .a(EX18), .b(EX20), .O(N1537) );
and2 gate227( .a(N614), .b(N957), .O(N1551) );
inv1 gate( .a(N1029),.O(N1029_NOT) );
inv1 gate( .a(N636),.O(N636_NOT));
and2 gate( .a(N1029_NOT), .b(p9), .O(EX21) );
and2 gate( .a(N636_NOT), .b(EX21), .O(EX22) );
and2 gate( .a(N1029), .b(p10), .O(EX23) );
and2 gate( .a(N636_NOT), .b(EX23), .O(EX24) );
and2 gate( .a(N1029_NOT), .b(p11), .O(EX25) );
and2 gate( .a(N636), .b(EX25), .O(EX26) );
and2 gate( .a(N1029), .b(p12), .O(EX27) );
and2 gate( .a(N636), .b(EX27), .O(EX28) );
or2  gate( .a(EX22), .b(EX24), .O(EX29) );
or2  gate( .a(EX26), .b(EX29), .O(EX30) );
or2  gate( .a(EX28), .b(EX30), .O(N1649) );
buf1 gate229( .a(N957), .O(N1703) );
nor2 gate230( .a(N957), .b(N614), .O(N1708) );
buf1 gate231( .a(N957), .O(N1713) );
nor2 gate232( .a(N614), .b(N957), .O(N1721) );
buf1 gate233( .a(N1029), .O(N1758) );
inv1 gate( .a(N163),.O(N163_NOT) );
inv1 gate( .a(N1116),.O(N1116_NOT));
and2 gate( .a(N163_NOT), .b(p13), .O(EX31) );
and2 gate( .a(N1116_NOT), .b(EX31), .O(EX32) );
and2 gate( .a(N163), .b(p14), .O(EX33) );
and2 gate( .a(N1116_NOT), .b(EX33), .O(EX34) );
and2 gate( .a(N163_NOT), .b(p15), .O(EX35) );
and2 gate( .a(N1116), .b(EX35), .O(EX36) );
and2 gate( .a(N163), .b(p16), .O(EX37) );
and2 gate( .a(N1116), .b(EX37), .O(EX38) );
or2  gate( .a(EX32), .b(EX34), .O(EX39) );
or2  gate( .a(EX36), .b(EX39), .O(EX40) );
or2  gate( .a(EX38), .b(EX40), .O(N1781) );
and2 gate235( .a(N170), .b(N1125), .O(N1782) );
inv1 gate236( .a(N1125), .O(N1783) );
inv1 gate237( .a(N1136), .O(N1789) );
and2 gate238( .a(N169), .b(N1125), .O(N1793) );
and2 gate239( .a(N168), .b(N1125), .O(N1794) );
and2 gate240( .a(N167), .b(N1125), .O(N1795) );
and2 gate241( .a(N166), .b(N1136), .O(N1796) );
and2 gate242( .a(N165), .b(N1136), .O(N1797) );
and2 gate243( .a(N164), .b(N1136), .O(N1798) );
inv1 gate244( .a(N1147), .O(N1799) );
inv1 gate245( .a(N1160), .O(N1805) );
and2 gate246( .a(N177), .b(N1147), .O(N1811) );
and2 gate247( .a(N176), .b(N1147), .O(N1812) );
and2 gate248( .a(N175), .b(N1147), .O(N1813) );
and2 gate249( .a(N174), .b(N1147), .O(N1814) );
and2 gate250( .a(N173), .b(N1147), .O(N1815) );
and2 gate251( .a(N157), .b(N1160), .O(N1816) );
and2 gate252( .a(N156), .b(N1160), .O(N1817) );
and2 gate253( .a(N155), .b(N1160), .O(N1818) );
and2 gate254( .a(N154), .b(N1160), .O(N1819) );
inv1 gate( .a(N153),.O(N153_NOT) );
inv1 gate( .a(N1160),.O(N1160_NOT));
and2 gate( .a(N153_NOT), .b(p17), .O(EX41) );
and2 gate( .a(N1160_NOT), .b(EX41), .O(EX42) );
and2 gate( .a(N153), .b(p18), .O(EX43) );
and2 gate( .a(N1160_NOT), .b(EX43), .O(EX44) );
and2 gate( .a(N153_NOT), .b(p19), .O(EX45) );
and2 gate( .a(N1160), .b(EX45), .O(EX46) );
and2 gate( .a(N153), .b(p20), .O(EX47) );
and2 gate( .a(N1160), .b(EX47), .O(EX48) );
or2  gate( .a(EX42), .b(EX44), .O(EX49) );
or2  gate( .a(EX46), .b(EX49), .O(EX50) );
or2  gate( .a(EX48), .b(EX50), .O(N1820) );
inv1 gate256( .a(N1284), .O(N1821) );
inv1 gate257( .a(N1287), .O(N1822) );
inv1 gate258( .a(N1290), .O(N1828) );
inv1 gate259( .a(N1293), .O(N1829) );
inv1 gate260( .a(N1296), .O(N1830) );
inv1 gate261( .a(N1299), .O(N1832) );
inv1 gate262( .a(N1302), .O(N1833) );
inv1 gate263( .a(N1305), .O(N1834) );
inv1 gate264( .a(N1308), .O(N1835) );
inv1 gate265( .a(N1311), .O(N1839) );
inv1 gate266( .a(N1314), .O(N1840) );
inv1 gate267( .a(N1317), .O(N1841) );
inv1 gate268( .a(N1320), .O(N1842) );
inv1 gate269( .a(N1323), .O(N1843) );
inv1 gate270( .a(N1175), .O(N1845) );
inv1 gate271( .a(N1182), .O(N1851) );
and2 gate272( .a(N181), .b(N1175), .O(N1857) );
and2 gate273( .a(N171), .b(N1175), .O(N1858) );
and2 gate274( .a(N180), .b(N1175), .O(N1859) );
and2 gate275( .a(N179), .b(N1175), .O(N1860) );
inv1 gate( .a(N178),.O(N178_NOT) );
inv1 gate( .a(N1175),.O(N1175_NOT));
and2 gate( .a(N178_NOT), .b(p21), .O(EX51) );
and2 gate( .a(N1175_NOT), .b(EX51), .O(EX52) );
and2 gate( .a(N178), .b(p22), .O(EX53) );
and2 gate( .a(N1175_NOT), .b(EX53), .O(EX54) );
and2 gate( .a(N178_NOT), .b(p23), .O(EX55) );
and2 gate( .a(N1175), .b(EX55), .O(EX56) );
and2 gate( .a(N178), .b(p24), .O(EX57) );
and2 gate( .a(N1175), .b(EX57), .O(EX58) );
or2  gate( .a(EX52), .b(EX54), .O(EX59) );
or2  gate( .a(EX56), .b(EX59), .O(EX60) );
or2  gate( .a(EX58), .b(EX60), .O(N1861) );
inv1 gate( .a(N161),.O(N161_NOT) );
inv1 gate( .a(N1182),.O(N1182_NOT));
and2 gate( .a(N161_NOT), .b(p25), .O(EX61) );
and2 gate( .a(N1182_NOT), .b(EX61), .O(EX62) );
and2 gate( .a(N161), .b(p26), .O(EX63) );
and2 gate( .a(N1182_NOT), .b(EX63), .O(EX64) );
and2 gate( .a(N161_NOT), .b(p27), .O(EX65) );
and2 gate( .a(N1182), .b(EX65), .O(EX66) );
and2 gate( .a(N161), .b(p28), .O(EX67) );
and2 gate( .a(N1182), .b(EX67), .O(EX68) );
or2  gate( .a(EX62), .b(EX64), .O(EX69) );
or2  gate( .a(EX66), .b(EX69), .O(EX70) );
or2  gate( .a(EX68), .b(EX70), .O(N1862) );
and2 gate278( .a(N151), .b(N1182), .O(N1863) );
and2 gate279( .a(N160), .b(N1182), .O(N1864) );
and2 gate280( .a(N159), .b(N1182), .O(N1865) );
and2 gate281( .a(N158), .b(N1182), .O(N1866) );
inv1 gate282( .a(N1326), .O(N1867) );
inv1 gate283( .a(N1329), .O(N1868) );
inv1 gate284( .a(N1332), .O(N1869) );
inv1 gate285( .a(N1335), .O(N1870) );
inv1 gate286( .a(N1338), .O(N1871) );
inv1 gate287( .a(N1341), .O(N1872) );
inv1 gate288( .a(N1344), .O(N1873) );
inv1 gate289( .a(N1347), .O(N1874) );
inv1 gate290( .a(N1350), .O(N1875) );
inv1 gate291( .a(N1353), .O(N1876) );
inv1 gate292( .a(N1356), .O(N1877) );
inv1 gate293( .a(N1359), .O(N1878) );
inv1 gate294( .a(N1362), .O(N1879) );
inv1 gate295( .a(N1365), .O(N1880) );
inv1 gate296( .a(N1368), .O(N1881) );
inv1 gate297( .a(N1371), .O(N1882) );
inv1 gate298( .a(N1374), .O(N1883) );
inv1 gate299( .a(N1377), .O(N1884) );
buf1 gate300( .a(N1199), .O(N1885) );
buf1 gate301( .a(N1194), .O(N1892) );
buf1 gate302( .a(N1199), .O(N1899) );
buf1 gate303( .a(N1194), .O(N1906) );
inv1 gate304( .a(N1211), .O(N1913) );
buf1 gate305( .a(N1194), .O(N1919) );
and2 gate306( .a(N44), .b(N1211), .O(N1926) );
and2 gate307( .a(N41), .b(N1211), .O(N1927) );
inv1 gate( .a(N29),.O(N29_NOT) );
inv1 gate( .a(N1211),.O(N1211_NOT));
and2 gate( .a(N29_NOT), .b(p29), .O(EX71) );
and2 gate( .a(N1211_NOT), .b(EX71), .O(EX72) );
and2 gate( .a(N29), .b(p30), .O(EX73) );
and2 gate( .a(N1211_NOT), .b(EX73), .O(EX74) );
and2 gate( .a(N29_NOT), .b(p31), .O(EX75) );
and2 gate( .a(N1211), .b(EX75), .O(EX76) );
and2 gate( .a(N29), .b(p32), .O(EX77) );
and2 gate( .a(N1211), .b(EX77), .O(EX78) );
or2  gate( .a(EX72), .b(EX74), .O(EX79) );
or2  gate( .a(EX76), .b(EX79), .O(EX80) );
or2  gate( .a(EX78), .b(EX80), .O(N1928) );
and2 gate309( .a(N26), .b(N1211), .O(N1929) );
and2 gate310( .a(N23), .b(N1211), .O(N1930) );
inv1 gate311( .a(N1380), .O(N1931) );
inv1 gate312( .a(N1383), .O(N1932) );
inv1 gate313( .a(N1386), .O(N1933) );
inv1 gate314( .a(N1389), .O(N1934) );
inv1 gate315( .a(N1392), .O(N1935) );
inv1 gate316( .a(N1395), .O(N1936) );
inv1 gate317( .a(N1398), .O(N1937) );
inv1 gate318( .a(N1401), .O(N1938) );
inv1 gate319( .a(N1404), .O(N1939) );
inv1 gate320( .a(N1407), .O(N1940) );
inv1 gate321( .a(N1410), .O(N1941) );
inv1 gate322( .a(N1413), .O(N1942) );
inv1 gate323( .a(N1416), .O(N1943) );
inv1 gate324( .a(N1419), .O(N1944) );
inv1 gate325( .a(N1422), .O(N1945) );
inv1 gate326( .a(N1425), .O(N1946) );
inv1 gate327( .a(N1233), .O(N1947) );
inv1 gate328( .a(N1244), .O(N1953) );
and2 gate329( .a(N209), .b(N1233), .O(N1957) );
and2 gate330( .a(N216), .b(N1233), .O(N1958) );
and2 gate331( .a(N215), .b(N1233), .O(N1959) );
and2 gate332( .a(N214), .b(N1233), .O(N1960) );
and2 gate333( .a(N213), .b(N1244), .O(N1961) );
and2 gate334( .a(N212), .b(N1244), .O(N1962) );
and2 gate335( .a(N211), .b(N1244), .O(N1963) );
inv1 gate336( .a(N1428), .O(N1965) );
and2 gate337( .a(N1222), .b(N636), .O(N1966) );
inv1 gate338( .a(N1431), .O(N1967) );
inv1 gate339( .a(N1434), .O(N1968) );
inv1 gate340( .a(N1437), .O(N1969) );
inv1 gate341( .a(N1440), .O(N1970) );
inv1 gate342( .a(N1443), .O(N1971) );
inv1 gate343( .a(N1446), .O(N1972) );
inv1 gate344( .a(N1449), .O(N1973) );
inv1 gate345( .a(N1452), .O(N1974) );
inv1 gate346( .a(N1455), .O(N1975) );
inv1 gate347( .a(N1458), .O(N1976) );
inv1 gate348( .a(N1249), .O(N1977) );
inv1 gate349( .a(N1256), .O(N1983) );
inv1 gate( .a(N642),.O(N642_NOT) );
inv1 gate( .a(N1249),.O(N1249_NOT));
and2 gate( .a(N642_NOT), .b(p33), .O(EX81) );
and2 gate( .a(N1249_NOT), .b(EX81), .O(EX82) );
and2 gate( .a(N642), .b(p34), .O(EX83) );
and2 gate( .a(N1249_NOT), .b(EX83), .O(EX84) );
and2 gate( .a(N642_NOT), .b(p35), .O(EX85) );
and2 gate( .a(N1249), .b(EX85), .O(EX86) );
and2 gate( .a(N642), .b(p36), .O(EX87) );
and2 gate( .a(N1249), .b(EX87), .O(EX88) );
or2  gate( .a(EX82), .b(EX84), .O(EX89) );
or2  gate( .a(EX86), .b(EX89), .O(EX90) );
or2  gate( .a(EX88), .b(EX90), .O(N1989) );
and2 gate351( .a(N644), .b(N1249), .O(N1990) );
and2 gate352( .a(N651), .b(N1249), .O(N1991) );
and2 gate353( .a(N674), .b(N1249), .O(N1992) );
and2 gate354( .a(N660), .b(N1249), .O(N1993) );
and2 gate355( .a(N666), .b(N1256), .O(N1994) );
and2 gate356( .a(N672), .b(N1256), .O(N1995) );
and2 gate357( .a(N673), .b(N1256), .O(N1996) );
inv1 gate358( .a(N1263), .O(N1997) );
buf1 gate359( .a(N1194), .O(N2003) );
and2 gate360( .a(N47), .b(N1263), .O(N2010) );
and2 gate361( .a(N35), .b(N1263), .O(N2011) );
and2 gate362( .a(N32), .b(N1263), .O(N2012) );
and2 gate363( .a(N50), .b(N1263), .O(N2013) );
and2 gate364( .a(N66), .b(N1263), .O(N2014) );
inv1 gate365( .a(N1461), .O(N2015) );
inv1 gate366( .a(N1464), .O(N2016) );
inv1 gate367( .a(N1467), .O(N2017) );
inv1 gate368( .a(N1470), .O(N2018) );
inv1 gate369( .a(N1473), .O(N2019) );
inv1 gate370( .a(N1476), .O(N2020) );
inv1 gate371( .a(N1479), .O(N2021) );
inv1 gate372( .a(N1482), .O(N2022) );
inv1 gate373( .a(N1485), .O(N2023) );
buf1 gate374( .a(N1206), .O(N2024) );
buf1 gate375( .a(N1206), .O(N2031) );
buf1 gate376( .a(N1206), .O(N2038) );
buf1 gate377( .a(N1206), .O(N2045) );
inv1 gate378( .a(N1270), .O(N2052) );
inv1 gate379( .a(N1277), .O(N2058) );
and2 gate380( .a(N706), .b(N1270), .O(N2064) );
and2 gate381( .a(N708), .b(N1270), .O(N2065) );
and2 gate382( .a(N715), .b(N1270), .O(N2066) );
inv1 gate( .a(N721),.O(N721_NOT) );
inv1 gate( .a(N1270),.O(N1270_NOT));
and2 gate( .a(N721_NOT), .b(p37), .O(EX91) );
and2 gate( .a(N1270_NOT), .b(EX91), .O(EX92) );
and2 gate( .a(N721), .b(p38), .O(EX93) );
and2 gate( .a(N1270_NOT), .b(EX93), .O(EX94) );
and2 gate( .a(N721_NOT), .b(p39), .O(EX95) );
and2 gate( .a(N1270), .b(EX95), .O(EX96) );
and2 gate( .a(N721), .b(p40), .O(EX97) );
and2 gate( .a(N1270), .b(EX97), .O(EX98) );
or2  gate( .a(EX92), .b(EX94), .O(EX99) );
or2  gate( .a(EX96), .b(EX99), .O(EX100) );
or2  gate( .a(EX98), .b(EX100), .O(N2067) );
inv1 gate( .a(N727),.O(N727_NOT) );
inv1 gate( .a(N1270),.O(N1270_NOT));
and2 gate( .a(N727_NOT), .b(p41), .O(EX101) );
and2 gate( .a(N1270_NOT), .b(EX101), .O(EX102) );
and2 gate( .a(N727), .b(p42), .O(EX103) );
and2 gate( .a(N1270_NOT), .b(EX103), .O(EX104) );
and2 gate( .a(N727_NOT), .b(p43), .O(EX105) );
and2 gate( .a(N1270), .b(EX105), .O(EX106) );
and2 gate( .a(N727), .b(p44), .O(EX107) );
and2 gate( .a(N1270), .b(EX107), .O(EX108) );
or2  gate( .a(EX102), .b(EX104), .O(EX109) );
or2  gate( .a(EX106), .b(EX109), .O(EX110) );
or2  gate( .a(EX108), .b(EX110), .O(N2068) );
and2 gate385( .a(N733), .b(N1277), .O(N2069) );
inv1 gate( .a(N734),.O(N734_NOT) );
inv1 gate( .a(N1277),.O(N1277_NOT));
and2 gate( .a(N734_NOT), .b(p45), .O(EX111) );
and2 gate( .a(N1277_NOT), .b(EX111), .O(EX112) );
and2 gate( .a(N734), .b(p46), .O(EX113) );
and2 gate( .a(N1277_NOT), .b(EX113), .O(EX114) );
and2 gate( .a(N734_NOT), .b(p47), .O(EX115) );
and2 gate( .a(N1277), .b(EX115), .O(EX116) );
and2 gate( .a(N734), .b(p48), .O(EX117) );
and2 gate( .a(N1277), .b(EX117), .O(EX118) );
or2  gate( .a(EX112), .b(EX114), .O(EX119) );
or2  gate( .a(EX116), .b(EX119), .O(EX120) );
or2  gate( .a(EX118), .b(EX120), .O(N2070) );
and2 gate387( .a(N742), .b(N1277), .O(N2071) );
and2 gate388( .a(N748), .b(N1277), .O(N2072) );
and2 gate389( .a(N749), .b(N1277), .O(N2073) );
buf1 gate390( .a(N1189), .O(N2074) );
buf1 gate391( .a(N1189), .O(N2081) );
buf1 gate392( .a(N1222), .O(N2086) );
nand2 gate393( .a(N1287), .b(N1821), .O(N2107) );
nand2 gate394( .a(N1284), .b(N1822), .O(N2108) );
inv1 gate395( .a(N1703), .O(N2110) );
nand2 gate396( .a(N1703), .b(N1832), .O(N2111) );
nand2 gate397( .a(N1308), .b(N1834), .O(N2112) );
nand2 gate398( .a(N1305), .b(N1835), .O(N2113) );
inv1 gate399( .a(N1713), .O(N2114) );
nand2 gate400( .a(N1713), .b(N1839), .O(N2115) );
inv1 gate401( .a(N1721), .O(N2117) );
inv1 gate402( .a(N1758), .O(N2171) );
nand2 gate403( .a(N1758), .b(N1965), .O(N2172) );
inv1 gate404( .a(N1708), .O(N2230) );
buf1 gate405( .a(N1537), .O(N2231) );
buf1 gate406( .a(N1551), .O(N2235) );
or2 gate407( .a(N1783), .b(N1782), .O(N2239) );
or2 gate408( .a(N1783), .b(N1125), .O(N2240) );
or2 gate409( .a(N1783), .b(N1793), .O(N2241) );
or2 gate410( .a(N1783), .b(N1794), .O(N2242) );
or2 gate411( .a(N1783), .b(N1795), .O(N2243) );
or2 gate412( .a(N1789), .b(N1796), .O(N2244) );
or2 gate413( .a(N1789), .b(N1797), .O(N2245) );
or2 gate414( .a(N1789), .b(N1798), .O(N2246) );
or2 gate415( .a(N1799), .b(N1811), .O(N2247) );
or2 gate416( .a(N1799), .b(N1812), .O(N2248) );
or2 gate417( .a(N1799), .b(N1813), .O(N2249) );
inv1 gate( .a(N1799),.O(N1799_NOT) );
inv1 gate( .a(N1814),.O(N1814_NOT));
and2 gate( .a(N1799_NOT), .b(p49), .O(EX121) );
and2 gate( .a(N1814_NOT), .b(EX121), .O(EX122) );
and2 gate( .a(N1799), .b(p50), .O(EX123) );
and2 gate( .a(N1814_NOT), .b(EX123), .O(EX124) );
and2 gate( .a(N1799_NOT), .b(p51), .O(EX125) );
and2 gate( .a(N1814), .b(EX125), .O(EX126) );
and2 gate( .a(N1799), .b(p52), .O(EX127) );
and2 gate( .a(N1814), .b(EX127), .O(EX128) );
or2  gate( .a(EX122), .b(EX124), .O(EX129) );
or2  gate( .a(EX126), .b(EX129), .O(EX130) );
or2  gate( .a(EX128), .b(EX130), .O(N2250) );
or2 gate419( .a(N1799), .b(N1815), .O(N2251) );
or2 gate420( .a(N1805), .b(N1816), .O(N2252) );
or2 gate421( .a(N1805), .b(N1817), .O(N2253) );
or2 gate422( .a(N1805), .b(N1818), .O(N2254) );
or2 gate423( .a(N1805), .b(N1819), .O(N2255) );
or2 gate424( .a(N1805), .b(N1820), .O(N2256) );
nand2 gate425( .a(N2107), .b(N2108), .O(N2257) );
inv1 gate426( .a(N2074), .O(N2267) );
nand2 gate427( .a(N1299), .b(N2110), .O(N2268) );
nand2 gate428( .a(N2112), .b(N2113), .O(N2269) );
nand2 gate429( .a(N1311), .b(N2114), .O(N2274) );
inv1 gate430( .a(N2081), .O(N2275) );
inv1 gate( .a(N141),.O(N141_NOT) );
inv1 gate( .a(N1845),.O(N1845_NOT));
and2 gate( .a(N141_NOT), .b(p53), .O(EX131) );
and2 gate( .a(N1845_NOT), .b(EX131), .O(EX132) );
and2 gate( .a(N141), .b(p54), .O(EX133) );
and2 gate( .a(N1845_NOT), .b(EX133), .O(EX134) );
and2 gate( .a(N141_NOT), .b(p55), .O(EX135) );
and2 gate( .a(N1845), .b(EX135), .O(EX136) );
and2 gate( .a(N141), .b(p56), .O(EX137) );
and2 gate( .a(N1845), .b(EX137), .O(EX138) );
or2  gate( .a(EX132), .b(EX134), .O(EX139) );
or2  gate( .a(EX136), .b(EX139), .O(EX140) );
or2  gate( .a(EX138), .b(EX140), .O(N2277) );
and2 gate432( .a(N147), .b(N1845), .O(N2278) );
inv1 gate( .a(N138),.O(N138_NOT) );
inv1 gate( .a(N1845),.O(N1845_NOT));
and2 gate( .a(N138_NOT), .b(p57), .O(EX141) );
and2 gate( .a(N1845_NOT), .b(EX141), .O(EX142) );
and2 gate( .a(N138), .b(p58), .O(EX143) );
and2 gate( .a(N1845_NOT), .b(EX143), .O(EX144) );
and2 gate( .a(N138_NOT), .b(p59), .O(EX145) );
and2 gate( .a(N1845), .b(EX145), .O(EX146) );
and2 gate( .a(N138), .b(p60), .O(EX147) );
and2 gate( .a(N1845), .b(EX147), .O(EX148) );
or2  gate( .a(EX142), .b(EX144), .O(EX149) );
or2  gate( .a(EX146), .b(EX149), .O(EX150) );
or2  gate( .a(EX148), .b(EX150), .O(N2279) );
and2 gate434( .a(N144), .b(N1845), .O(N2280) );
inv1 gate( .a(N135),.O(N135_NOT) );
inv1 gate( .a(N1845),.O(N1845_NOT));
and2 gate( .a(N135_NOT), .b(p61), .O(EX151) );
and2 gate( .a(N1845_NOT), .b(EX151), .O(EX152) );
and2 gate( .a(N135), .b(p62), .O(EX153) );
and2 gate( .a(N1845_NOT), .b(EX153), .O(EX154) );
and2 gate( .a(N135_NOT), .b(p63), .O(EX155) );
and2 gate( .a(N1845), .b(EX155), .O(EX156) );
and2 gate( .a(N135), .b(p64), .O(EX157) );
and2 gate( .a(N1845), .b(EX157), .O(EX158) );
or2  gate( .a(EX152), .b(EX154), .O(EX159) );
or2  gate( .a(EX156), .b(EX159), .O(EX160) );
or2  gate( .a(EX158), .b(EX160), .O(N2281) );
inv1 gate( .a(N141),.O(N141_NOT) );
inv1 gate( .a(N1851),.O(N1851_NOT));
and2 gate( .a(N141_NOT), .b(p65), .O(EX161) );
and2 gate( .a(N1851_NOT), .b(EX161), .O(EX162) );
and2 gate( .a(N141), .b(p66), .O(EX163) );
and2 gate( .a(N1851_NOT), .b(EX163), .O(EX164) );
and2 gate( .a(N141_NOT), .b(p67), .O(EX165) );
and2 gate( .a(N1851), .b(EX165), .O(EX166) );
and2 gate( .a(N141), .b(p68), .O(EX167) );
and2 gate( .a(N1851), .b(EX167), .O(EX168) );
or2  gate( .a(EX162), .b(EX164), .O(EX169) );
or2  gate( .a(EX166), .b(EX169), .O(EX170) );
or2  gate( .a(EX168), .b(EX170), .O(N2282) );
and2 gate437( .a(N147), .b(N1851), .O(N2283) );
and2 gate438( .a(N138), .b(N1851), .O(N2284) );
and2 gate439( .a(N144), .b(N1851), .O(N2285) );
inv1 gate( .a(N135),.O(N135_NOT) );
inv1 gate( .a(N1851),.O(N1851_NOT));
and2 gate( .a(N135_NOT), .b(p69), .O(EX171) );
and2 gate( .a(N1851_NOT), .b(EX171), .O(EX172) );
and2 gate( .a(N135), .b(p70), .O(EX173) );
and2 gate( .a(N1851_NOT), .b(EX173), .O(EX174) );
and2 gate( .a(N135_NOT), .b(p71), .O(EX175) );
and2 gate( .a(N1851), .b(EX175), .O(EX176) );
and2 gate( .a(N135), .b(p72), .O(EX177) );
and2 gate( .a(N1851), .b(EX177), .O(EX178) );
or2  gate( .a(EX172), .b(EX174), .O(EX179) );
or2  gate( .a(EX176), .b(EX179), .O(EX180) );
or2  gate( .a(EX178), .b(EX180), .O(N2286) );
inv1 gate441( .a(N1885), .O(N2287) );
inv1 gate442( .a(N1892), .O(N2293) );
and2 gate443( .a(N103), .b(N1885), .O(N2299) );
and2 gate444( .a(N130), .b(N1885), .O(N2300) );
and2 gate445( .a(N127), .b(N1885), .O(N2301) );
inv1 gate( .a(N124),.O(N124_NOT) );
inv1 gate( .a(N1885),.O(N1885_NOT));
and2 gate( .a(N124_NOT), .b(p73), .O(EX181) );
and2 gate( .a(N1885_NOT), .b(EX181), .O(EX182) );
and2 gate( .a(N124), .b(p74), .O(EX183) );
and2 gate( .a(N1885_NOT), .b(EX183), .O(EX184) );
and2 gate( .a(N124_NOT), .b(p75), .O(EX185) );
and2 gate( .a(N1885), .b(EX185), .O(EX186) );
and2 gate( .a(N124), .b(p76), .O(EX187) );
and2 gate( .a(N1885), .b(EX187), .O(EX188) );
or2  gate( .a(EX182), .b(EX184), .O(EX189) );
or2  gate( .a(EX186), .b(EX189), .O(EX190) );
or2  gate( .a(EX188), .b(EX190), .O(N2302) );
and2 gate447( .a(N100), .b(N1885), .O(N2303) );
inv1 gate( .a(N103),.O(N103_NOT) );
inv1 gate( .a(N1892),.O(N1892_NOT));
and2 gate( .a(N103_NOT), .b(p77), .O(EX191) );
and2 gate( .a(N1892_NOT), .b(EX191), .O(EX192) );
and2 gate( .a(N103), .b(p78), .O(EX193) );
and2 gate( .a(N1892_NOT), .b(EX193), .O(EX194) );
and2 gate( .a(N103_NOT), .b(p79), .O(EX195) );
and2 gate( .a(N1892), .b(EX195), .O(EX196) );
and2 gate( .a(N103), .b(p80), .O(EX197) );
and2 gate( .a(N1892), .b(EX197), .O(EX198) );
or2  gate( .a(EX192), .b(EX194), .O(EX199) );
or2  gate( .a(EX196), .b(EX199), .O(EX200) );
or2  gate( .a(EX198), .b(EX200), .O(N2304) );
and2 gate449( .a(N130), .b(N1892), .O(N2305) );
and2 gate450( .a(N127), .b(N1892), .O(N2306) );
and2 gate451( .a(N124), .b(N1892), .O(N2307) );
and2 gate452( .a(N100), .b(N1892), .O(N2308) );
inv1 gate453( .a(N1899), .O(N2309) );
inv1 gate454( .a(N1906), .O(N2315) );
inv1 gate( .a(N115),.O(N115_NOT) );
inv1 gate( .a(N1899),.O(N1899_NOT));
and2 gate( .a(N115_NOT), .b(p81), .O(EX201) );
and2 gate( .a(N1899_NOT), .b(EX201), .O(EX202) );
and2 gate( .a(N115), .b(p82), .O(EX203) );
and2 gate( .a(N1899_NOT), .b(EX203), .O(EX204) );
and2 gate( .a(N115_NOT), .b(p83), .O(EX205) );
and2 gate( .a(N1899), .b(EX205), .O(EX206) );
and2 gate( .a(N115), .b(p84), .O(EX207) );
and2 gate( .a(N1899), .b(EX207), .O(EX208) );
or2  gate( .a(EX202), .b(EX204), .O(EX209) );
or2  gate( .a(EX206), .b(EX209), .O(EX210) );
or2  gate( .a(EX208), .b(EX210), .O(N2321) );
and2 gate456( .a(N118), .b(N1899), .O(N2322) );
and2 gate457( .a(N97), .b(N1899), .O(N2323) );
and2 gate458( .a(N94), .b(N1899), .O(N2324) );
and2 gate459( .a(N121), .b(N1899), .O(N2325) );
and2 gate460( .a(N115), .b(N1906), .O(N2326) );
and2 gate461( .a(N118), .b(N1906), .O(N2327) );
and2 gate462( .a(N97), .b(N1906), .O(N2328) );
and2 gate463( .a(N94), .b(N1906), .O(N2329) );
and2 gate464( .a(N121), .b(N1906), .O(N2330) );
inv1 gate465( .a(N1919), .O(N2331) );
and2 gate466( .a(N208), .b(N1913), .O(N2337) );
and2 gate467( .a(N198), .b(N1913), .O(N2338) );
and2 gate468( .a(N207), .b(N1913), .O(N2339) );
and2 gate469( .a(N206), .b(N1913), .O(N2340) );
and2 gate470( .a(N205), .b(N1913), .O(N2341) );
and2 gate471( .a(N44), .b(N1919), .O(N2342) );
inv1 gate( .a(N41),.O(N41_NOT) );
inv1 gate( .a(N1919),.O(N1919_NOT));
and2 gate( .a(N41_NOT), .b(p85), .O(EX211) );
and2 gate( .a(N1919_NOT), .b(EX211), .O(EX212) );
and2 gate( .a(N41), .b(p86), .O(EX213) );
and2 gate( .a(N1919_NOT), .b(EX213), .O(EX214) );
and2 gate( .a(N41_NOT), .b(p87), .O(EX215) );
and2 gate( .a(N1919), .b(EX215), .O(EX216) );
and2 gate( .a(N41), .b(p88), .O(EX217) );
and2 gate( .a(N1919), .b(EX217), .O(EX218) );
or2  gate( .a(EX212), .b(EX214), .O(EX219) );
or2  gate( .a(EX216), .b(EX219), .O(EX220) );
or2  gate( .a(EX218), .b(EX220), .O(N2343) );
and2 gate473( .a(N29), .b(N1919), .O(N2344) );
and2 gate474( .a(N26), .b(N1919), .O(N2345) );
and2 gate475( .a(N23), .b(N1919), .O(N2346) );
inv1 gate( .a(N1947),.O(N1947_NOT) );
inv1 gate( .a(N1233),.O(N1233_NOT));
and2 gate( .a(N1947_NOT), .b(p89), .O(EX221) );
and2 gate( .a(N1233_NOT), .b(EX221), .O(EX222) );
and2 gate( .a(N1947), .b(p90), .O(EX223) );
and2 gate( .a(N1233_NOT), .b(EX223), .O(EX224) );
and2 gate( .a(N1947_NOT), .b(p91), .O(EX225) );
and2 gate( .a(N1233), .b(EX225), .O(EX226) );
and2 gate( .a(N1947), .b(p92), .O(EX227) );
and2 gate( .a(N1233), .b(EX227), .O(EX228) );
or2  gate( .a(EX222), .b(EX224), .O(EX229) );
or2  gate( .a(EX226), .b(EX229), .O(EX230) );
or2  gate( .a(EX228), .b(EX230), .O(N2347) );
or2 gate477( .a(N1947), .b(N1957), .O(N2348) );
or2 gate478( .a(N1947), .b(N1958), .O(N2349) );
or2 gate479( .a(N1947), .b(N1959), .O(N2350) );
or2 gate480( .a(N1947), .b(N1960), .O(N2351) );
or2 gate481( .a(N1953), .b(N1961), .O(N2352) );
or2 gate482( .a(N1953), .b(N1962), .O(N2353) );
or2 gate483( .a(N1953), .b(N1963), .O(N2354) );
nand2 gate484( .a(N1428), .b(N2171), .O(N2355) );
inv1 gate485( .a(N2086), .O(N2356) );
nand2 gate486( .a(N2086), .b(N1967), .O(N2357) );
and2 gate487( .a(N114), .b(N1977), .O(N2358) );
and2 gate488( .a(N113), .b(N1977), .O(N2359) );
and2 gate489( .a(N111), .b(N1977), .O(N2360) );
and2 gate490( .a(N87), .b(N1977), .O(N2361) );
and2 gate491( .a(N112), .b(N1977), .O(N2362) );
and2 gate492( .a(N88), .b(N1983), .O(N2363) );
and2 gate493( .a(N245), .b(N1983), .O(N2364) );
and2 gate494( .a(N271), .b(N1983), .O(N2365) );
and2 gate495( .a(N759), .b(N1983), .O(N2366) );
and2 gate496( .a(N70), .b(N1983), .O(N2367) );
inv1 gate497( .a(N2003), .O(N2368) );
and2 gate498( .a(N193), .b(N1997), .O(N2374) );
and2 gate499( .a(N192), .b(N1997), .O(N2375) );
and2 gate500( .a(N191), .b(N1997), .O(N2376) );
and2 gate501( .a(N190), .b(N1997), .O(N2377) );
and2 gate502( .a(N189), .b(N1997), .O(N2378) );
and2 gate503( .a(N47), .b(N2003), .O(N2379) );
and2 gate504( .a(N35), .b(N2003), .O(N2380) );
and2 gate505( .a(N32), .b(N2003), .O(N2381) );
and2 gate506( .a(N50), .b(N2003), .O(N2382) );
and2 gate507( .a(N66), .b(N2003), .O(N2383) );
inv1 gate508( .a(N2024), .O(N2384) );
inv1 gate509( .a(N2031), .O(N2390) );
and2 gate510( .a(N58), .b(N2024), .O(N2396) );
inv1 gate( .a(N77),.O(N77_NOT) );
inv1 gate( .a(N2024),.O(N2024_NOT));
and2 gate( .a(N77_NOT), .b(p93), .O(EX231) );
and2 gate( .a(N2024_NOT), .b(EX231), .O(EX232) );
and2 gate( .a(N77), .b(p94), .O(EX233) );
and2 gate( .a(N2024_NOT), .b(EX233), .O(EX234) );
and2 gate( .a(N77_NOT), .b(p95), .O(EX235) );
and2 gate( .a(N2024), .b(EX235), .O(EX236) );
and2 gate( .a(N77), .b(p96), .O(EX237) );
and2 gate( .a(N2024), .b(EX237), .O(EX238) );
or2  gate( .a(EX232), .b(EX234), .O(EX239) );
or2  gate( .a(EX236), .b(EX239), .O(EX240) );
or2  gate( .a(EX238), .b(EX240), .O(N2397) );
and2 gate512( .a(N78), .b(N2024), .O(N2398) );
and2 gate513( .a(N59), .b(N2024), .O(N2399) );
and2 gate514( .a(N81), .b(N2024), .O(N2400) );
and2 gate515( .a(N80), .b(N2031), .O(N2401) );
inv1 gate( .a(N79),.O(N79_NOT) );
inv1 gate( .a(N2031),.O(N2031_NOT));
and2 gate( .a(N79_NOT), .b(p97), .O(EX241) );
and2 gate( .a(N2031_NOT), .b(EX241), .O(EX242) );
and2 gate( .a(N79), .b(p98), .O(EX243) );
and2 gate( .a(N2031_NOT), .b(EX243), .O(EX244) );
and2 gate( .a(N79_NOT), .b(p99), .O(EX245) );
and2 gate( .a(N2031), .b(EX245), .O(EX246) );
and2 gate( .a(N79), .b(p100), .O(EX247) );
and2 gate( .a(N2031), .b(EX247), .O(EX248) );
or2  gate( .a(EX242), .b(EX244), .O(EX249) );
or2  gate( .a(EX246), .b(EX249), .O(EX250) );
or2  gate( .a(EX248), .b(EX250), .O(N2402) );
and2 gate517( .a(N60), .b(N2031), .O(N2403) );
and2 gate518( .a(N61), .b(N2031), .O(N2404) );
and2 gate519( .a(N62), .b(N2031), .O(N2405) );
inv1 gate520( .a(N2038), .O(N2406) );
inv1 gate521( .a(N2045), .O(N2412) );
and2 gate522( .a(N69), .b(N2038), .O(N2418) );
and2 gate523( .a(N70), .b(N2038), .O(N2419) );
and2 gate524( .a(N74), .b(N2038), .O(N2420) );
and2 gate525( .a(N76), .b(N2038), .O(N2421) );
and2 gate526( .a(N75), .b(N2038), .O(N2422) );
and2 gate527( .a(N73), .b(N2045), .O(N2423) );
and2 gate528( .a(N53), .b(N2045), .O(N2424) );
and2 gate529( .a(N54), .b(N2045), .O(N2425) );
and2 gate530( .a(N55), .b(N2045), .O(N2426) );
and2 gate531( .a(N56), .b(N2045), .O(N2427) );
and2 gate532( .a(N82), .b(N2052), .O(N2428) );
and2 gate533( .a(N65), .b(N2052), .O(N2429) );
and2 gate534( .a(N83), .b(N2052), .O(N2430) );
inv1 gate( .a(N84),.O(N84_NOT) );
inv1 gate( .a(N2052),.O(N2052_NOT));
and2 gate( .a(N84_NOT), .b(p101), .O(EX251) );
and2 gate( .a(N2052_NOT), .b(EX251), .O(EX252) );
and2 gate( .a(N84), .b(p102), .O(EX253) );
and2 gate( .a(N2052_NOT), .b(EX253), .O(EX254) );
and2 gate( .a(N84_NOT), .b(p103), .O(EX255) );
and2 gate( .a(N2052), .b(EX255), .O(EX256) );
and2 gate( .a(N84), .b(p104), .O(EX257) );
and2 gate( .a(N2052), .b(EX257), .O(EX258) );
or2  gate( .a(EX252), .b(EX254), .O(EX259) );
or2  gate( .a(EX256), .b(EX259), .O(EX260) );
or2  gate( .a(EX258), .b(EX260), .O(N2431) );
and2 gate536( .a(N85), .b(N2052), .O(N2432) );
and2 gate537( .a(N64), .b(N2058), .O(N2433) );
and2 gate538( .a(N63), .b(N2058), .O(N2434) );
and2 gate539( .a(N86), .b(N2058), .O(N2435) );
inv1 gate( .a(N109),.O(N109_NOT) );
inv1 gate( .a(N2058),.O(N2058_NOT));
and2 gate( .a(N109_NOT), .b(p105), .O(EX261) );
and2 gate( .a(N2058_NOT), .b(EX261), .O(EX262) );
and2 gate( .a(N109), .b(p106), .O(EX263) );
and2 gate( .a(N2058_NOT), .b(EX263), .O(EX264) );
and2 gate( .a(N109_NOT), .b(p107), .O(EX265) );
and2 gate( .a(N2058), .b(EX265), .O(EX266) );
and2 gate( .a(N109), .b(p108), .O(EX267) );
and2 gate( .a(N2058), .b(EX267), .O(EX268) );
or2  gate( .a(EX262), .b(EX264), .O(EX269) );
or2  gate( .a(EX266), .b(EX269), .O(EX270) );
or2  gate( .a(EX268), .b(EX270), .O(N2436) );
and2 gate541( .a(N110), .b(N2058), .O(N2437) );
inv1 gate( .a(N2239),.O(N2239_NOT) );
inv1 gate( .a(N1119),.O(N1119_NOT));
and2 gate( .a(N2239_NOT), .b(p109), .O(EX271) );
and2 gate( .a(N1119_NOT), .b(EX271), .O(EX272) );
and2 gate( .a(N2239), .b(p110), .O(EX273) );
and2 gate( .a(N1119_NOT), .b(EX273), .O(EX274) );
and2 gate( .a(N2239_NOT), .b(p111), .O(EX275) );
and2 gate( .a(N1119), .b(EX275), .O(EX276) );
and2 gate( .a(N2239), .b(p112), .O(EX277) );
and2 gate( .a(N1119), .b(EX277), .O(EX278) );
or2  gate( .a(EX272), .b(EX274), .O(EX279) );
or2  gate( .a(EX276), .b(EX279), .O(EX280) );
or2  gate( .a(EX278), .b(EX280), .O(N2441) );
and2 gate543( .a(N2240), .b(N1119), .O(N2442) );
and2 gate544( .a(N2241), .b(N1119), .O(N2446) );
inv1 gate( .a(N2242),.O(N2242_NOT) );
inv1 gate( .a(N1119),.O(N1119_NOT));
and2 gate( .a(N2242_NOT), .b(p113), .O(EX281) );
and2 gate( .a(N1119_NOT), .b(EX281), .O(EX282) );
and2 gate( .a(N2242), .b(p114), .O(EX283) );
and2 gate( .a(N1119_NOT), .b(EX283), .O(EX284) );
and2 gate( .a(N2242_NOT), .b(p115), .O(EX285) );
and2 gate( .a(N1119), .b(EX285), .O(EX286) );
and2 gate( .a(N2242), .b(p116), .O(EX287) );
and2 gate( .a(N1119), .b(EX287), .O(EX288) );
or2  gate( .a(EX282), .b(EX284), .O(EX289) );
or2  gate( .a(EX286), .b(EX289), .O(EX290) );
or2  gate( .a(EX288), .b(EX290), .O(N2450) );
and2 gate546( .a(N2243), .b(N1119), .O(N2454) );
and2 gate547( .a(N2244), .b(N1132), .O(N2458) );
and2 gate548( .a(N2247), .b(N1141), .O(N2462) );
and2 gate549( .a(N2248), .b(N1141), .O(N2466) );
and2 gate550( .a(N2249), .b(N1141), .O(N2470) );
inv1 gate( .a(N2250),.O(N2250_NOT) );
inv1 gate( .a(N1141),.O(N1141_NOT));
and2 gate( .a(N2250_NOT), .b(p117), .O(EX291) );
and2 gate( .a(N1141_NOT), .b(EX291), .O(EX292) );
and2 gate( .a(N2250), .b(p118), .O(EX293) );
and2 gate( .a(N1141_NOT), .b(EX293), .O(EX294) );
and2 gate( .a(N2250_NOT), .b(p119), .O(EX295) );
and2 gate( .a(N1141), .b(EX295), .O(EX296) );
and2 gate( .a(N2250), .b(p120), .O(EX297) );
and2 gate( .a(N1141), .b(EX297), .O(EX298) );
or2  gate( .a(EX292), .b(EX294), .O(EX299) );
or2  gate( .a(EX296), .b(EX299), .O(EX300) );
or2  gate( .a(EX298), .b(EX300), .O(N2474) );
and2 gate552( .a(N2251), .b(N1141), .O(N2478) );
and2 gate553( .a(N2252), .b(N1154), .O(N2482) );
and2 gate554( .a(N2253), .b(N1154), .O(N2488) );
and2 gate555( .a(N2254), .b(N1154), .O(N2496) );
and2 gate556( .a(N2255), .b(N1154), .O(N2502) );
and2 gate557( .a(N2256), .b(N1154), .O(N2508) );
nand2 gate558( .a(N2268), .b(N2111), .O(N2523) );
nand2 gate559( .a(N2274), .b(N2115), .O(N2533) );
inv1 gate560( .a(N2235), .O(N2537) );
or2 gate561( .a(N2278), .b(N1858), .O(N2538) );
or2 gate562( .a(N2279), .b(N1859), .O(N2542) );
or2 gate563( .a(N2280), .b(N1860), .O(N2546) );
or2 gate564( .a(N2281), .b(N1861), .O(N2550) );
or2 gate565( .a(N2283), .b(N1863), .O(N2554) );
or2 gate566( .a(N2284), .b(N1864), .O(N2561) );
or2 gate567( .a(N2285), .b(N1865), .O(N2567) );
or2 gate568( .a(N2286), .b(N1866), .O(N2573) );
or2 gate569( .a(N2338), .b(N1927), .O(N2604) );
or2 gate570( .a(N2339), .b(N1928), .O(N2607) );
inv1 gate( .a(N2340),.O(N2340_NOT) );
inv1 gate( .a(N1929),.O(N1929_NOT));
and2 gate( .a(N2340_NOT), .b(p121), .O(EX301) );
and2 gate( .a(N1929_NOT), .b(EX301), .O(EX302) );
and2 gate( .a(N2340), .b(p122), .O(EX303) );
and2 gate( .a(N1929_NOT), .b(EX303), .O(EX304) );
and2 gate( .a(N2340_NOT), .b(p123), .O(EX305) );
and2 gate( .a(N1929), .b(EX305), .O(EX306) );
and2 gate( .a(N2340), .b(p124), .O(EX307) );
and2 gate( .a(N1929), .b(EX307), .O(EX308) );
or2  gate( .a(EX302), .b(EX304), .O(EX309) );
or2  gate( .a(EX306), .b(EX309), .O(EX310) );
or2  gate( .a(EX308), .b(EX310), .O(N2611) );
or2 gate572( .a(N2341), .b(N1930), .O(N2615) );
and2 gate573( .a(N2348), .b(N1227), .O(N2619) );
inv1 gate( .a(N2349),.O(N2349_NOT) );
inv1 gate( .a(N1227),.O(N1227_NOT));
and2 gate( .a(N2349_NOT), .b(p125), .O(EX311) );
and2 gate( .a(N1227_NOT), .b(EX311), .O(EX312) );
and2 gate( .a(N2349), .b(p126), .O(EX313) );
and2 gate( .a(N1227_NOT), .b(EX313), .O(EX314) );
and2 gate( .a(N2349_NOT), .b(p127), .O(EX315) );
and2 gate( .a(N1227), .b(EX315), .O(EX316) );
and2 gate( .a(N2349), .b(p128), .O(EX317) );
and2 gate( .a(N1227), .b(EX317), .O(EX318) );
or2  gate( .a(EX312), .b(EX314), .O(EX319) );
or2  gate( .a(EX316), .b(EX319), .O(EX320) );
or2  gate( .a(EX318), .b(EX320), .O(N2626) );
and2 gate575( .a(N2350), .b(N1227), .O(N2632) );
and2 gate576( .a(N2351), .b(N1227), .O(N2638) );
and2 gate577( .a(N2352), .b(N1240), .O(N2644) );
inv1 gate( .a(N2355),.O(N2355_NOT) );
inv1 gate( .a(N2172),.O(N2172_NOT));
and2 gate( .a(N2355_NOT), .b(p129), .O(EX321) );
and2 gate( .a(N2172_NOT), .b(EX321), .O(EX322) );
and2 gate( .a(N2355), .b(p130), .O(EX323) );
and2 gate( .a(N2172_NOT), .b(EX323), .O(EX324) );
and2 gate( .a(N2355_NOT), .b(p131), .O(EX325) );
and2 gate( .a(N2172), .b(EX325), .O(EX326) );
and2 gate( .a(N2355), .b(p132), .O(EX327) );
and2 gate( .a(N2172), .b(EX327), .O(EX328) );
or2  gate( .a(EX322), .b(EX324), .O(EX329) );
or2  gate( .a(EX326), .b(EX329), .O(EX330) );
or2  gate( .a(EX328), .b(EX330), .O(N2650) );
nand2 gate579( .a(N1431), .b(N2356), .O(N2653) );
or2 gate580( .a(N2359), .b(N1990), .O(N2654) );
or2 gate581( .a(N2360), .b(N1991), .O(N2658) );
or2 gate582( .a(N2361), .b(N1992), .O(N2662) );
or2 gate583( .a(N2362), .b(N1993), .O(N2666) );
or2 gate584( .a(N2363), .b(N1994), .O(N2670) );
or2 gate585( .a(N2366), .b(N1256), .O(N2674) );
inv1 gate( .a(N2367),.O(N2367_NOT) );
inv1 gate( .a(N1256),.O(N1256_NOT));
and2 gate( .a(N2367_NOT), .b(p133), .O(EX331) );
and2 gate( .a(N1256_NOT), .b(EX331), .O(EX332) );
and2 gate( .a(N2367), .b(p134), .O(EX333) );
and2 gate( .a(N1256_NOT), .b(EX333), .O(EX334) );
and2 gate( .a(N2367_NOT), .b(p135), .O(EX335) );
and2 gate( .a(N1256), .b(EX335), .O(EX336) );
and2 gate( .a(N2367), .b(p136), .O(EX337) );
and2 gate( .a(N1256), .b(EX337), .O(EX338) );
or2  gate( .a(EX332), .b(EX334), .O(EX339) );
or2  gate( .a(EX336), .b(EX339), .O(EX340) );
or2  gate( .a(EX338), .b(EX340), .O(N2680) );
or2 gate587( .a(N2374), .b(N2010), .O(N2688) );
or2 gate588( .a(N2375), .b(N2011), .O(N2692) );
or2 gate589( .a(N2376), .b(N2012), .O(N2696) );
or2 gate590( .a(N2377), .b(N2013), .O(N2700) );
or2 gate591( .a(N2378), .b(N2014), .O(N2704) );
and2 gate592( .a(N2347), .b(N1227), .O(N2728) );
or2 gate593( .a(N2429), .b(N2065), .O(N2729) );
or2 gate594( .a(N2430), .b(N2066), .O(N2733) );
or2 gate595( .a(N2431), .b(N2067), .O(N2737) );
or2 gate596( .a(N2432), .b(N2068), .O(N2741) );
or2 gate597( .a(N2433), .b(N2069), .O(N2745) );
or2 gate598( .a(N2434), .b(N2070), .O(N2749) );
or2 gate599( .a(N2435), .b(N2071), .O(N2753) );
inv1 gate( .a(N2436),.O(N2436_NOT) );
inv1 gate( .a(N2072),.O(N2072_NOT));
and2 gate( .a(N2436_NOT), .b(p137), .O(EX341) );
and2 gate( .a(N2072_NOT), .b(EX341), .O(EX342) );
and2 gate( .a(N2436), .b(p138), .O(EX343) );
and2 gate( .a(N2072_NOT), .b(EX343), .O(EX344) );
and2 gate( .a(N2436_NOT), .b(p139), .O(EX345) );
and2 gate( .a(N2072), .b(EX345), .O(EX346) );
and2 gate( .a(N2436), .b(p140), .O(EX347) );
and2 gate( .a(N2072), .b(EX347), .O(EX348) );
or2  gate( .a(EX342), .b(EX344), .O(EX349) );
or2  gate( .a(EX346), .b(EX349), .O(EX350) );
or2  gate( .a(EX348), .b(EX350), .O(N2757) );
or2 gate601( .a(N2437), .b(N2073), .O(N2761) );
inv1 gate602( .a(N2231), .O(N2765) );
inv1 gate( .a(N2354),.O(N2354_NOT) );
inv1 gate( .a(N1240),.O(N1240_NOT));
and2 gate( .a(N2354_NOT), .b(p141), .O(EX351) );
and2 gate( .a(N1240_NOT), .b(EX351), .O(EX352) );
and2 gate( .a(N2354), .b(p142), .O(EX353) );
and2 gate( .a(N1240_NOT), .b(EX353), .O(EX354) );
and2 gate( .a(N2354_NOT), .b(p143), .O(EX355) );
and2 gate( .a(N1240), .b(EX355), .O(EX356) );
and2 gate( .a(N2354), .b(p144), .O(EX357) );
and2 gate( .a(N1240), .b(EX357), .O(EX358) );
or2  gate( .a(EX352), .b(EX354), .O(EX359) );
or2  gate( .a(EX356), .b(EX359), .O(EX360) );
or2  gate( .a(EX358), .b(EX360), .O(N2766) );
and2 gate604( .a(N2353), .b(N1240), .O(N2769) );
and2 gate605( .a(N2246), .b(N1132), .O(N2772) );
and2 gate606( .a(N2245), .b(N1132), .O(N2775) );
or2 gate607( .a(N2282), .b(N1862), .O(N2778) );
inv1 gate( .a(N2358),.O(N2358_NOT) );
inv1 gate( .a(N1989),.O(N1989_NOT));
and2 gate( .a(N2358_NOT), .b(p145), .O(EX361) );
and2 gate( .a(N1989_NOT), .b(EX361), .O(EX362) );
and2 gate( .a(N2358), .b(p146), .O(EX363) );
and2 gate( .a(N1989_NOT), .b(EX363), .O(EX364) );
and2 gate( .a(N2358_NOT), .b(p147), .O(EX365) );
and2 gate( .a(N1989), .b(EX365), .O(EX366) );
and2 gate( .a(N2358), .b(p148), .O(EX367) );
and2 gate( .a(N1989), .b(EX367), .O(EX368) );
or2  gate( .a(EX362), .b(EX364), .O(EX369) );
or2  gate( .a(EX366), .b(EX369), .O(EX370) );
or2  gate( .a(EX368), .b(EX370), .O(N2781) );
inv1 gate( .a(N2365),.O(N2365_NOT) );
inv1 gate( .a(N1996),.O(N1996_NOT));
and2 gate( .a(N2365_NOT), .b(p149), .O(EX371) );
and2 gate( .a(N1996_NOT), .b(EX371), .O(EX372) );
and2 gate( .a(N2365), .b(p150), .O(EX373) );
and2 gate( .a(N1996_NOT), .b(EX373), .O(EX374) );
and2 gate( .a(N2365_NOT), .b(p151), .O(EX375) );
and2 gate( .a(N1996), .b(EX375), .O(EX376) );
and2 gate( .a(N2365), .b(p152), .O(EX377) );
and2 gate( .a(N1996), .b(EX377), .O(EX378) );
or2  gate( .a(EX372), .b(EX374), .O(EX379) );
or2  gate( .a(EX376), .b(EX379), .O(EX380) );
or2  gate( .a(EX378), .b(EX380), .O(N2784) );
or2 gate610( .a(N2364), .b(N1995), .O(N2787) );
or2 gate611( .a(N2337), .b(N1926), .O(N2790) );
or2 gate612( .a(N2277), .b(N1857), .O(N2793) );
or2 gate613( .a(N2428), .b(N2064), .O(N2796) );
inv1 gate( .a(N2257),.O(N2257_NOT) );
inv1 gate( .a(N1537),.O(N1537_NOT));
and2 gate( .a(N2257_NOT), .b(p153), .O(EX381) );
and2 gate( .a(N1537_NOT), .b(EX381), .O(EX382) );
and2 gate( .a(N2257), .b(p154), .O(EX383) );
and2 gate( .a(N1537_NOT), .b(EX383), .O(EX384) );
and2 gate( .a(N2257_NOT), .b(p155), .O(EX385) );
and2 gate( .a(N1537), .b(EX385), .O(EX386) );
and2 gate( .a(N2257), .b(p156), .O(EX387) );
and2 gate( .a(N1537), .b(EX387), .O(EX388) );
or2  gate( .a(EX382), .b(EX384), .O(EX389) );
or2  gate( .a(EX386), .b(EX389), .O(EX390) );
or2  gate( .a(EX388), .b(EX390), .O(N2866) );
and2 gate615( .a(N2257), .b(N1537), .O(N2867) );
and2 gate616( .a(N2257), .b(N1537), .O(N2868) );
and2 gate617( .a(N2257), .b(N1537), .O(N2869) );
and2 gate618( .a(N2269), .b(N1551), .O(N2878) );
and2 gate619( .a(N204), .b(N2287), .O(N2913) );
and2 gate620( .a(N203), .b(N2287), .O(N2914) );
inv1 gate( .a(N202),.O(N202_NOT) );
inv1 gate( .a(N2287),.O(N2287_NOT));
and2 gate( .a(N202_NOT), .b(p157), .O(EX391) );
and2 gate( .a(N2287_NOT), .b(EX391), .O(EX392) );
and2 gate( .a(N202), .b(p158), .O(EX393) );
and2 gate( .a(N2287_NOT), .b(EX393), .O(EX394) );
and2 gate( .a(N202_NOT), .b(p159), .O(EX395) );
and2 gate( .a(N2287), .b(EX395), .O(EX396) );
and2 gate( .a(N202), .b(p160), .O(EX397) );
and2 gate( .a(N2287), .b(EX397), .O(EX398) );
or2  gate( .a(EX392), .b(EX394), .O(EX399) );
or2  gate( .a(EX396), .b(EX399), .O(EX400) );
or2  gate( .a(EX398), .b(EX400), .O(N2915) );
and2 gate622( .a(N201), .b(N2287), .O(N2916) );
and2 gate623( .a(N200), .b(N2287), .O(N2917) );
and2 gate624( .a(N235), .b(N2293), .O(N2918) );
and2 gate625( .a(N234), .b(N2293), .O(N2919) );
and2 gate626( .a(N233), .b(N2293), .O(N2920) );
and2 gate627( .a(N232), .b(N2293), .O(N2921) );
and2 gate628( .a(N231), .b(N2293), .O(N2922) );
and2 gate629( .a(N197), .b(N2309), .O(N2923) );
and2 gate630( .a(N187), .b(N2309), .O(N2924) );
and2 gate631( .a(N196), .b(N2309), .O(N2925) );
and2 gate632( .a(N195), .b(N2309), .O(N2926) );
and2 gate633( .a(N194), .b(N2309), .O(N2927) );
and2 gate634( .a(N227), .b(N2315), .O(N2928) );
and2 gate635( .a(N217), .b(N2315), .O(N2929) );
and2 gate636( .a(N226), .b(N2315), .O(N2930) );
and2 gate637( .a(N225), .b(N2315), .O(N2931) );
and2 gate638( .a(N224), .b(N2315), .O(N2932) );
and2 gate639( .a(N239), .b(N2331), .O(N2933) );
and2 gate640( .a(N229), .b(N2331), .O(N2934) );
and2 gate641( .a(N238), .b(N2331), .O(N2935) );
and2 gate642( .a(N237), .b(N2331), .O(N2936) );
and2 gate643( .a(N236), .b(N2331), .O(N2937) );
nand2 gate644( .a(N2653), .b(N2357), .O(N2988) );
and2 gate645( .a(N223), .b(N2368), .O(N3005) );
and2 gate646( .a(N222), .b(N2368), .O(N3006) );
and2 gate647( .a(N221), .b(N2368), .O(N3007) );
and2 gate648( .a(N220), .b(N2368), .O(N3008) );
and2 gate649( .a(N219), .b(N2368), .O(N3009) );
and2 gate650( .a(N812), .b(N2384), .O(N3020) );
and2 gate651( .a(N814), .b(N2384), .O(N3021) );
inv1 gate( .a(N821),.O(N821_NOT) );
inv1 gate( .a(N2384),.O(N2384_NOT));
and2 gate( .a(N821_NOT), .b(p161), .O(EX401) );
and2 gate( .a(N2384_NOT), .b(EX401), .O(EX402) );
and2 gate( .a(N821), .b(p162), .O(EX403) );
and2 gate( .a(N2384_NOT), .b(EX403), .O(EX404) );
and2 gate( .a(N821_NOT), .b(p163), .O(EX405) );
and2 gate( .a(N2384), .b(EX405), .O(EX406) );
and2 gate( .a(N821), .b(p164), .O(EX407) );
and2 gate( .a(N2384), .b(EX407), .O(EX408) );
or2  gate( .a(EX402), .b(EX404), .O(EX409) );
or2  gate( .a(EX406), .b(EX409), .O(EX410) );
or2  gate( .a(EX408), .b(EX410), .O(N3022) );
and2 gate653( .a(N827), .b(N2384), .O(N3023) );
and2 gate654( .a(N833), .b(N2384), .O(N3024) );
and2 gate655( .a(N839), .b(N2390), .O(N3025) );
and2 gate656( .a(N845), .b(N2390), .O(N3026) );
and2 gate657( .a(N853), .b(N2390), .O(N3027) );
and2 gate658( .a(N859), .b(N2390), .O(N3028) );
and2 gate659( .a(N865), .b(N2390), .O(N3029) );
and2 gate660( .a(N758), .b(N2406), .O(N3032) );
and2 gate661( .a(N759), .b(N2406), .O(N3033) );
and2 gate662( .a(N762), .b(N2406), .O(N3034) );
and2 gate663( .a(N768), .b(N2406), .O(N3035) );
and2 gate664( .a(N774), .b(N2406), .O(N3036) );
and2 gate665( .a(N780), .b(N2412), .O(N3037) );
and2 gate666( .a(N786), .b(N2412), .O(N3038) );
and2 gate667( .a(N794), .b(N2412), .O(N3039) );
and2 gate668( .a(N800), .b(N2412), .O(N3040) );
and2 gate669( .a(N806), .b(N2412), .O(N3041) );
buf1 gate670( .a(N2257), .O(N3061) );
buf1 gate671( .a(N2257), .O(N3064) );
buf1 gate672( .a(N2269), .O(N3067) );
buf1 gate673( .a(N2269), .O(N3070) );
inv1 gate674( .a(N2728), .O(N3073) );
inv1 gate675( .a(N2441), .O(N3080) );
inv1 gate( .a(N666),.O(N666_NOT) );
inv1 gate( .a(N2644),.O(N2644_NOT));
and2 gate( .a(N666_NOT), .b(p165), .O(EX411) );
and2 gate( .a(N2644_NOT), .b(EX411), .O(EX412) );
and2 gate( .a(N666), .b(p166), .O(EX413) );
and2 gate( .a(N2644_NOT), .b(EX413), .O(EX414) );
and2 gate( .a(N666_NOT), .b(p167), .O(EX415) );
and2 gate( .a(N2644), .b(EX415), .O(EX416) );
and2 gate( .a(N666), .b(p168), .O(EX417) );
and2 gate( .a(N2644), .b(EX417), .O(EX418) );
or2  gate( .a(EX412), .b(EX414), .O(EX419) );
or2  gate( .a(EX416), .b(EX419), .O(EX420) );
or2  gate( .a(EX418), .b(EX420), .O(N3096) );
and2 gate677( .a(N660), .b(N2638), .O(N3097) );
and2 gate678( .a(N1189), .b(N2632), .O(N3101) );
and2 gate679( .a(N651), .b(N2626), .O(N3107) );
and2 gate680( .a(N644), .b(N2619), .O(N3114) );
and2 gate681( .a(N2523), .b(N2257), .O(N3122) );
inv1 gate( .a(N1167),.O(N1167_NOT) );
inv1 gate( .a(N2866),.O(N2866_NOT));
and2 gate( .a(N1167_NOT), .b(p169), .O(EX421) );
and2 gate( .a(N2866_NOT), .b(EX421), .O(EX422) );
and2 gate( .a(N1167), .b(p170), .O(EX423) );
and2 gate( .a(N2866_NOT), .b(EX423), .O(EX424) );
and2 gate( .a(N1167_NOT), .b(p171), .O(EX425) );
and2 gate( .a(N2866), .b(EX425), .O(EX426) );
and2 gate( .a(N1167), .b(p172), .O(EX427) );
and2 gate( .a(N2866), .b(EX427), .O(EX428) );
or2  gate( .a(EX422), .b(EX424), .O(EX429) );
or2  gate( .a(EX426), .b(EX429), .O(EX430) );
or2  gate( .a(EX428), .b(EX430), .O(N3126) );
and2 gate683( .a(N2523), .b(N2257), .O(N3130) );
or2 gate684( .a(N1167), .b(N2869), .O(N3131) );
and2 gate685( .a(N2523), .b(N2257), .O(N3134) );
inv1 gate686( .a(N2533), .O(N3135) );
and2 gate687( .a(N666), .b(N2644), .O(N3136) );
inv1 gate( .a(N660),.O(N660_NOT) );
inv1 gate( .a(N2638),.O(N2638_NOT));
and2 gate( .a(N660_NOT), .b(p173), .O(EX431) );
and2 gate( .a(N2638_NOT), .b(EX431), .O(EX432) );
and2 gate( .a(N660), .b(p174), .O(EX433) );
and2 gate( .a(N2638_NOT), .b(EX433), .O(EX434) );
and2 gate( .a(N660_NOT), .b(p175), .O(EX435) );
and2 gate( .a(N2638), .b(EX435), .O(EX436) );
and2 gate( .a(N660), .b(p176), .O(EX437) );
and2 gate( .a(N2638), .b(EX437), .O(EX438) );
or2  gate( .a(EX432), .b(EX434), .O(EX439) );
or2  gate( .a(EX436), .b(EX439), .O(EX440) );
or2  gate( .a(EX438), .b(EX440), .O(N3137) );
and2 gate689( .a(N1189), .b(N2632), .O(N3140) );
inv1 gate( .a(N651),.O(N651_NOT) );
inv1 gate( .a(N2626),.O(N2626_NOT));
and2 gate( .a(N651_NOT), .b(p177), .O(EX441) );
and2 gate( .a(N2626_NOT), .b(EX441), .O(EX442) );
and2 gate( .a(N651), .b(p178), .O(EX443) );
and2 gate( .a(N2626_NOT), .b(EX443), .O(EX444) );
and2 gate( .a(N651_NOT), .b(p179), .O(EX445) );
and2 gate( .a(N2626), .b(EX445), .O(EX446) );
and2 gate( .a(N651), .b(p180), .O(EX447) );
and2 gate( .a(N2626), .b(EX447), .O(EX448) );
or2  gate( .a(EX442), .b(EX444), .O(EX449) );
or2  gate( .a(EX446), .b(EX449), .O(EX450) );
or2  gate( .a(EX448), .b(EX450), .O(N3144) );
and2 gate691( .a(N644), .b(N2619), .O(N3149) );
and2 gate692( .a(N2533), .b(N2269), .O(N3155) );
or2 gate693( .a(N1174), .b(N2878), .O(N3159) );
inv1 gate694( .a(N2778), .O(N3167) );
and2 gate695( .a(N609), .b(N2508), .O(N3168) );
and2 gate696( .a(N604), .b(N2502), .O(N3169) );
and2 gate697( .a(N742), .b(N2496), .O(N3173) );
and2 gate698( .a(N734), .b(N2488), .O(N3178) );
and2 gate699( .a(N599), .b(N2482), .O(N3184) );
and2 gate700( .a(N727), .b(N2573), .O(N3185) );
and2 gate701( .a(N721), .b(N2567), .O(N3189) );
and2 gate702( .a(N715), .b(N2561), .O(N3195) );
and2 gate703( .a(N708), .b(N2554), .O(N3202) );
and2 gate704( .a(N609), .b(N2508), .O(N3210) );
and2 gate705( .a(N604), .b(N2502), .O(N3211) );
and2 gate706( .a(N742), .b(N2496), .O(N3215) );
and2 gate707( .a(N2488), .b(N734), .O(N3221) );
inv1 gate( .a(N599),.O(N599_NOT) );
inv1 gate( .a(N2482),.O(N2482_NOT));
and2 gate( .a(N599_NOT), .b(p181), .O(EX451) );
and2 gate( .a(N2482_NOT), .b(EX451), .O(EX452) );
and2 gate( .a(N599), .b(p182), .O(EX453) );
and2 gate( .a(N2482_NOT), .b(EX453), .O(EX454) );
and2 gate( .a(N599_NOT), .b(p183), .O(EX455) );
and2 gate( .a(N2482), .b(EX455), .O(EX456) );
and2 gate( .a(N599), .b(p184), .O(EX457) );
and2 gate( .a(N2482), .b(EX457), .O(EX458) );
or2  gate( .a(EX452), .b(EX454), .O(EX459) );
or2  gate( .a(EX456), .b(EX459), .O(EX460) );
or2  gate( .a(EX458), .b(EX460), .O(N3228) );
and2 gate709( .a(N727), .b(N2573), .O(N3229) );
and2 gate710( .a(N721), .b(N2567), .O(N3232) );
inv1 gate( .a(N715),.O(N715_NOT) );
inv1 gate( .a(N2561),.O(N2561_NOT));
and2 gate( .a(N715_NOT), .b(p185), .O(EX461) );
and2 gate( .a(N2561_NOT), .b(EX461), .O(EX462) );
and2 gate( .a(N715), .b(p186), .O(EX463) );
and2 gate( .a(N2561_NOT), .b(EX463), .O(EX464) );
and2 gate( .a(N715_NOT), .b(p187), .O(EX465) );
and2 gate( .a(N2561), .b(EX465), .O(EX466) );
and2 gate( .a(N715), .b(p188), .O(EX467) );
and2 gate( .a(N2561), .b(EX467), .O(EX468) );
or2  gate( .a(EX462), .b(EX464), .O(EX469) );
or2  gate( .a(EX466), .b(EX469), .O(EX470) );
or2  gate( .a(EX468), .b(EX470), .O(N3236) );
and2 gate712( .a(N708), .b(N2554), .O(N3241) );
or2 gate713( .a(N2913), .b(N2299), .O(N3247) );
or2 gate714( .a(N2914), .b(N2300), .O(N3251) );
or2 gate715( .a(N2915), .b(N2301), .O(N3255) );
or2 gate716( .a(N2916), .b(N2302), .O(N3259) );
or2 gate717( .a(N2917), .b(N2303), .O(N3263) );
inv1 gate( .a(N2918),.O(N2918_NOT) );
inv1 gate( .a(N2304),.O(N2304_NOT));
and2 gate( .a(N2918_NOT), .b(p189), .O(EX471) );
and2 gate( .a(N2304_NOT), .b(EX471), .O(EX472) );
and2 gate( .a(N2918), .b(p190), .O(EX473) );
and2 gate( .a(N2304_NOT), .b(EX473), .O(EX474) );
and2 gate( .a(N2918_NOT), .b(p191), .O(EX475) );
and2 gate( .a(N2304), .b(EX475), .O(EX476) );
and2 gate( .a(N2918), .b(p192), .O(EX477) );
and2 gate( .a(N2304), .b(EX477), .O(EX478) );
or2  gate( .a(EX472), .b(EX474), .O(EX479) );
or2  gate( .a(EX476), .b(EX479), .O(EX480) );
or2  gate( .a(EX478), .b(EX480), .O(N3267) );
or2 gate719( .a(N2919), .b(N2305), .O(N3273) );
or2 gate720( .a(N2920), .b(N2306), .O(N3281) );
or2 gate721( .a(N2921), .b(N2307), .O(N3287) );
or2 gate722( .a(N2922), .b(N2308), .O(N3293) );
or2 gate723( .a(N2924), .b(N2322), .O(N3299) );
or2 gate724( .a(N2925), .b(N2323), .O(N3303) );
inv1 gate( .a(N2926),.O(N2926_NOT) );
inv1 gate( .a(N2324),.O(N2324_NOT));
and2 gate( .a(N2926_NOT), .b(p193), .O(EX481) );
and2 gate( .a(N2324_NOT), .b(EX481), .O(EX482) );
and2 gate( .a(N2926), .b(p194), .O(EX483) );
and2 gate( .a(N2324_NOT), .b(EX483), .O(EX484) );
and2 gate( .a(N2926_NOT), .b(p195), .O(EX485) );
and2 gate( .a(N2324), .b(EX485), .O(EX486) );
and2 gate( .a(N2926), .b(p196), .O(EX487) );
and2 gate( .a(N2324), .b(EX487), .O(EX488) );
or2  gate( .a(EX482), .b(EX484), .O(EX489) );
or2  gate( .a(EX486), .b(EX489), .O(EX490) );
or2  gate( .a(EX488), .b(EX490), .O(N3307) );
or2 gate726( .a(N2927), .b(N2325), .O(N3311) );
or2 gate727( .a(N2929), .b(N2327), .O(N3315) );
or2 gate728( .a(N2930), .b(N2328), .O(N3322) );
or2 gate729( .a(N2931), .b(N2329), .O(N3328) );
or2 gate730( .a(N2932), .b(N2330), .O(N3334) );
or2 gate731( .a(N2934), .b(N2343), .O(N3340) );
or2 gate732( .a(N2935), .b(N2344), .O(N3343) );
or2 gate733( .a(N2936), .b(N2345), .O(N3349) );
or2 gate734( .a(N2937), .b(N2346), .O(N3355) );
and2 gate735( .a(N2761), .b(N2478), .O(N3361) );
and2 gate736( .a(N2757), .b(N2474), .O(N3362) );
and2 gate737( .a(N2753), .b(N2470), .O(N3363) );
and2 gate738( .a(N2749), .b(N2466), .O(N3364) );
and2 gate739( .a(N2745), .b(N2462), .O(N3365) );
and2 gate740( .a(N2741), .b(N2550), .O(N3366) );
and2 gate741( .a(N2737), .b(N2546), .O(N3367) );
inv1 gate( .a(N2733),.O(N2733_NOT) );
inv1 gate( .a(N2542),.O(N2542_NOT));
and2 gate( .a(N2733_NOT), .b(p197), .O(EX491) );
and2 gate( .a(N2542_NOT), .b(EX491), .O(EX492) );
and2 gate( .a(N2733), .b(p198), .O(EX493) );
and2 gate( .a(N2542_NOT), .b(EX493), .O(EX494) );
and2 gate( .a(N2733_NOT), .b(p199), .O(EX495) );
and2 gate( .a(N2542), .b(EX495), .O(EX496) );
and2 gate( .a(N2733), .b(p200), .O(EX497) );
and2 gate( .a(N2542), .b(EX497), .O(EX498) );
or2  gate( .a(EX492), .b(EX494), .O(EX499) );
or2  gate( .a(EX496), .b(EX499), .O(EX500) );
or2  gate( .a(EX498), .b(EX500), .O(N3368) );
and2 gate743( .a(N2729), .b(N2538), .O(N3369) );
and2 gate744( .a(N2670), .b(N2458), .O(N3370) );
and2 gate745( .a(N2666), .b(N2454), .O(N3371) );
and2 gate746( .a(N2662), .b(N2450), .O(N3372) );
inv1 gate( .a(N2658),.O(N2658_NOT) );
inv1 gate( .a(N2446),.O(N2446_NOT));
and2 gate( .a(N2658_NOT), .b(p201), .O(EX501) );
and2 gate( .a(N2446_NOT), .b(EX501), .O(EX502) );
and2 gate( .a(N2658), .b(p202), .O(EX503) );
and2 gate( .a(N2446_NOT), .b(EX503), .O(EX504) );
and2 gate( .a(N2658_NOT), .b(p203), .O(EX505) );
and2 gate( .a(N2446), .b(EX505), .O(EX506) );
and2 gate( .a(N2658), .b(p204), .O(EX507) );
and2 gate( .a(N2446), .b(EX507), .O(EX508) );
or2  gate( .a(EX502), .b(EX504), .O(EX509) );
or2  gate( .a(EX506), .b(EX509), .O(EX510) );
or2  gate( .a(EX508), .b(EX510), .O(N3373) );
and2 gate748( .a(N2654), .b(N2442), .O(N3374) );
and2 gate749( .a(N2988), .b(N2650), .O(N3375) );
and2 gate750( .a(N2650), .b(N1966), .O(N3379) );
inv1 gate751( .a(N2781), .O(N3380) );
and2 gate752( .a(N695), .b(N2604), .O(N3381) );
or2 gate753( .a(N3005), .b(N2379), .O(N3384) );
or2 gate754( .a(N3006), .b(N2380), .O(N3390) );
or2 gate755( .a(N3007), .b(N2381), .O(N3398) );
or2 gate756( .a(N3008), .b(N2382), .O(N3404) );
or2 gate757( .a(N3009), .b(N2383), .O(N3410) );
or2 gate758( .a(N3021), .b(N2397), .O(N3416) );
or2 gate759( .a(N3022), .b(N2398), .O(N3420) );
or2 gate760( .a(N3023), .b(N2399), .O(N3424) );
or2 gate761( .a(N3024), .b(N2400), .O(N3428) );
or2 gate762( .a(N3025), .b(N2401), .O(N3432) );
or2 gate763( .a(N3026), .b(N2402), .O(N3436) );
or2 gate764( .a(N3027), .b(N2403), .O(N3440) );
or2 gate765( .a(N3028), .b(N2404), .O(N3444) );
or2 gate766( .a(N3029), .b(N2405), .O(N3448) );
inv1 gate767( .a(N2790), .O(N3452) );
inv1 gate768( .a(N2793), .O(N3453) );
or2 gate769( .a(N3034), .b(N2420), .O(N3454) );
or2 gate770( .a(N3035), .b(N2421), .O(N3458) );
or2 gate771( .a(N3036), .b(N2422), .O(N3462) );
or2 gate772( .a(N3037), .b(N2423), .O(N3466) );
or2 gate773( .a(N3038), .b(N2424), .O(N3470) );
or2 gate774( .a(N3039), .b(N2425), .O(N3474) );
or2 gate775( .a(N3040), .b(N2426), .O(N3478) );
or2 gate776( .a(N3041), .b(N2427), .O(N3482) );
inv1 gate777( .a(N2796), .O(N3486) );
buf1 gate778( .a(N2644), .O(N3487) );
buf1 gate779( .a(N2638), .O(N3490) );
buf1 gate780( .a(N2632), .O(N3493) );
buf1 gate781( .a(N2626), .O(N3496) );
buf1 gate782( .a(N2619), .O(N3499) );
buf1 gate783( .a(N2523), .O(N3502) );
nor2 gate784( .a(N1167), .b(N2868), .O(N3507) );
buf1 gate785( .a(N2523), .O(N3510) );
nor2 gate786( .a(N644), .b(N2619), .O(N3515) );
buf1 gate787( .a(N2644), .O(N3518) );
buf1 gate788( .a(N2638), .O(N3521) );
buf1 gate789( .a(N2632), .O(N3524) );
buf1 gate790( .a(N2626), .O(N3527) );
buf1 gate791( .a(N2619), .O(N3530) );
buf1 gate792( .a(N2619), .O(N3535) );
buf1 gate793( .a(N2632), .O(N3539) );
buf1 gate794( .a(N2626), .O(N3542) );
buf1 gate795( .a(N2644), .O(N3545) );
buf1 gate796( .a(N2638), .O(N3548) );
inv1 gate797( .a(N2766), .O(N3551) );
inv1 gate798( .a(N2769), .O(N3552) );
buf1 gate799( .a(N2442), .O(N3553) );
buf1 gate800( .a(N2450), .O(N3557) );
buf1 gate801( .a(N2446), .O(N3560) );
buf1 gate802( .a(N2458), .O(N3563) );
buf1 gate803( .a(N2454), .O(N3566) );
inv1 gate804( .a(N2772), .O(N3569) );
inv1 gate805( .a(N2775), .O(N3570) );
buf1 gate806( .a(N2554), .O(N3571) );
buf1 gate807( .a(N2567), .O(N3574) );
buf1 gate808( .a(N2561), .O(N3577) );
buf1 gate809( .a(N2482), .O(N3580) );
buf1 gate810( .a(N2573), .O(N3583) );
buf1 gate811( .a(N2496), .O(N3586) );
buf1 gate812( .a(N2488), .O(N3589) );
buf1 gate813( .a(N2508), .O(N3592) );
buf1 gate814( .a(N2502), .O(N3595) );
buf1 gate815( .a(N2508), .O(N3598) );
buf1 gate816( .a(N2502), .O(N3601) );
buf1 gate817( .a(N2496), .O(N3604) );
buf1 gate818( .a(N2482), .O(N3607) );
buf1 gate819( .a(N2573), .O(N3610) );
buf1 gate820( .a(N2567), .O(N3613) );
buf1 gate821( .a(N2561), .O(N3616) );
buf1 gate822( .a(N2488), .O(N3619) );
buf1 gate823( .a(N2554), .O(N3622) );
nor2 gate824( .a(N734), .b(N2488), .O(N3625) );
nor2 gate825( .a(N708), .b(N2554), .O(N3628) );
buf1 gate826( .a(N2508), .O(N3631) );
buf1 gate827( .a(N2502), .O(N3634) );
buf1 gate828( .a(N2496), .O(N3637) );
buf1 gate829( .a(N2488), .O(N3640) );
buf1 gate830( .a(N2482), .O(N3643) );
buf1 gate831( .a(N2573), .O(N3646) );
buf1 gate832( .a(N2567), .O(N3649) );
buf1 gate833( .a(N2561), .O(N3652) );
buf1 gate834( .a(N2554), .O(N3655) );
inv1 gate( .a(N2488),.O(N2488_NOT) );
inv1 gate( .a(N734),.O(N734_NOT));
and2 gate( .a(N2488_NOT), .b(p205), .O(EX511) );
and2 gate( .a(N734_NOT), .b(EX511), .O(EX512) );
and2 gate( .a(N2488), .b(p206), .O(EX513) );
and2 gate( .a(N734_NOT), .b(EX513), .O(EX514) );
and2 gate( .a(N2488_NOT), .b(p207), .O(EX515) );
and2 gate( .a(N734), .b(EX515), .O(EX516) );
and2 gate( .a(N2488), .b(p208), .O(EX517) );
and2 gate( .a(N734), .b(EX517), .O(EX518) );
or2  gate( .a(EX512), .b(EX514), .O(EX519) );
or2  gate( .a(EX516), .b(EX519), .O(EX520) );
or2  gate( .a(EX518), .b(EX520), .O(N3658) );
buf1 gate836( .a(N2674), .O(N3661) );
buf1 gate837( .a(N2674), .O(N3664) );
buf1 gate838( .a(N2761), .O(N3667) );
buf1 gate839( .a(N2478), .O(N3670) );
buf1 gate840( .a(N2757), .O(N3673) );
buf1 gate841( .a(N2474), .O(N3676) );
buf1 gate842( .a(N2753), .O(N3679) );
buf1 gate843( .a(N2470), .O(N3682) );
buf1 gate844( .a(N2745), .O(N3685) );
buf1 gate845( .a(N2462), .O(N3688) );
buf1 gate846( .a(N2741), .O(N3691) );
buf1 gate847( .a(N2550), .O(N3694) );
buf1 gate848( .a(N2737), .O(N3697) );
buf1 gate849( .a(N2546), .O(N3700) );
buf1 gate850( .a(N2733), .O(N3703) );
buf1 gate851( .a(N2542), .O(N3706) );
buf1 gate852( .a(N2749), .O(N3709) );
buf1 gate853( .a(N2466), .O(N3712) );
buf1 gate854( .a(N2729), .O(N3715) );
buf1 gate855( .a(N2538), .O(N3718) );
buf1 gate856( .a(N2704), .O(N3721) );
buf1 gate857( .a(N2700), .O(N3724) );
buf1 gate858( .a(N2696), .O(N3727) );
buf1 gate859( .a(N2688), .O(N3730) );
buf1 gate860( .a(N2692), .O(N3733) );
buf1 gate861( .a(N2670), .O(N3736) );
buf1 gate862( .a(N2458), .O(N3739) );
buf1 gate863( .a(N2666), .O(N3742) );
buf1 gate864( .a(N2454), .O(N3745) );
buf1 gate865( .a(N2662), .O(N3748) );
buf1 gate866( .a(N2450), .O(N3751) );
buf1 gate867( .a(N2658), .O(N3754) );
buf1 gate868( .a(N2446), .O(N3757) );
buf1 gate869( .a(N2654), .O(N3760) );
buf1 gate870( .a(N2442), .O(N3763) );
buf1 gate871( .a(N2654), .O(N3766) );
buf1 gate872( .a(N2662), .O(N3769) );
buf1 gate873( .a(N2658), .O(N3772) );
buf1 gate874( .a(N2670), .O(N3775) );
buf1 gate875( .a(N2666), .O(N3778) );
inv1 gate876( .a(N2784), .O(N3781) );
inv1 gate877( .a(N2787), .O(N3782) );
or2 gate878( .a(N2928), .b(N2326), .O(N3783) );
or2 gate879( .a(N2933), .b(N2342), .O(N3786) );
or2 gate880( .a(N2923), .b(N2321), .O(N3789) );
buf1 gate881( .a(N2688), .O(N3792) );
buf1 gate882( .a(N2696), .O(N3795) );
buf1 gate883( .a(N2692), .O(N3798) );
buf1 gate884( .a(N2704), .O(N3801) );
buf1 gate885( .a(N2700), .O(N3804) );
buf1 gate886( .a(N2604), .O(N3807) );
buf1 gate887( .a(N2611), .O(N3810) );
buf1 gate888( .a(N2607), .O(N3813) );
buf1 gate889( .a(N2615), .O(N3816) );
buf1 gate890( .a(N2538), .O(N3819) );
buf1 gate891( .a(N2546), .O(N3822) );
buf1 gate892( .a(N2542), .O(N3825) );
buf1 gate893( .a(N2462), .O(N3828) );
buf1 gate894( .a(N2550), .O(N3831) );
buf1 gate895( .a(N2470), .O(N3834) );
buf1 gate896( .a(N2466), .O(N3837) );
buf1 gate897( .a(N2478), .O(N3840) );
buf1 gate898( .a(N2474), .O(N3843) );
buf1 gate899( .a(N2615), .O(N3846) );
buf1 gate900( .a(N2611), .O(N3849) );
buf1 gate901( .a(N2607), .O(N3852) );
buf1 gate902( .a(N2680), .O(N3855) );
buf1 gate903( .a(N2729), .O(N3858) );
buf1 gate904( .a(N2737), .O(N3861) );
buf1 gate905( .a(N2733), .O(N3864) );
buf1 gate906( .a(N2745), .O(N3867) );
buf1 gate907( .a(N2741), .O(N3870) );
buf1 gate908( .a(N2753), .O(N3873) );
buf1 gate909( .a(N2749), .O(N3876) );
buf1 gate910( .a(N2761), .O(N3879) );
buf1 gate911( .a(N2757), .O(N3882) );
or2 gate912( .a(N3033), .b(N2419), .O(N3885) );
or2 gate913( .a(N3032), .b(N2418), .O(N3888) );
or2 gate914( .a(N3020), .b(N2396), .O(N3891) );
nand2 gate915( .a(N3067), .b(N2117), .O(N3953) );
inv1 gate916( .a(N3067), .O(N3954) );
inv1 gate( .a(N3070),.O(N3070_NOT) );
inv1 gate( .a(N2537),.O(N2537_NOT));
and2 gate( .a(N3070_NOT), .b(p209), .O(EX521) );
and2 gate( .a(N2537_NOT), .b(EX521), .O(EX522) );
and2 gate( .a(N3070), .b(p210), .O(EX523) );
and2 gate( .a(N2537_NOT), .b(EX523), .O(EX524) );
and2 gate( .a(N3070_NOT), .b(p211), .O(EX525) );
and2 gate( .a(N2537), .b(EX525), .O(EX526) );
and2 gate( .a(N3070), .b(p212), .O(EX527) );
and2 gate( .a(N2537), .b(EX527), .O(EX528) );
or2  gate( .a(EX522), .b(EX524), .O(EX529) );
or2  gate( .a(EX526), .b(EX529), .O(EX530) );
or2  gate( .a(EX528), .b(EX530), .O(N3955) );
inv1 gate918( .a(N3070), .O(N3956) );
inv1 gate919( .a(N3073), .O(N3958) );
inv1 gate920( .a(N3080), .O(N3964) );
or2 gate921( .a(N1649), .b(N3379), .O(N4193) );
or3 gate922( .a(N1167), .b(N2867), .c(N3130), .O(N4303) );
inv1 gate923( .a(N3061), .O(N4308) );
inv1 gate924( .a(N3064), .O(N4313) );
nand2 gate925( .a(N2769), .b(N3551), .O(N4326) );
nand2 gate926( .a(N2766), .b(N3552), .O(N4327) );
inv1 gate( .a(N2775),.O(N2775_NOT) );
inv1 gate( .a(N3569),.O(N3569_NOT));
and2 gate( .a(N2775_NOT), .b(p213), .O(EX531) );
and2 gate( .a(N3569_NOT), .b(EX531), .O(EX532) );
and2 gate( .a(N2775), .b(p214), .O(EX533) );
and2 gate( .a(N3569_NOT), .b(EX533), .O(EX534) );
and2 gate( .a(N2775_NOT), .b(p215), .O(EX535) );
and2 gate( .a(N3569), .b(EX535), .O(EX536) );
and2 gate( .a(N2775), .b(p216), .O(EX537) );
and2 gate( .a(N3569), .b(EX537), .O(EX538) );
or2  gate( .a(EX532), .b(EX534), .O(EX539) );
or2  gate( .a(EX536), .b(EX539), .O(EX540) );
or2  gate( .a(EX538), .b(EX540), .O(N4333) );
nand2 gate928( .a(N2772), .b(N3570), .O(N4334) );
nand2 gate929( .a(N2787), .b(N3781), .O(N4411) );
nand2 gate930( .a(N2784), .b(N3782), .O(N4412) );
nand2 gate931( .a(N3487), .b(N1828), .O(N4463) );
inv1 gate932( .a(N3487), .O(N4464) );
nand2 gate933( .a(N3490), .b(N1829), .O(N4465) );
inv1 gate934( .a(N3490), .O(N4466) );
nand2 gate935( .a(N3493), .b(N2267), .O(N4467) );
inv1 gate936( .a(N3493), .O(N4468) );
inv1 gate( .a(N3496),.O(N3496_NOT) );
inv1 gate( .a(N1830),.O(N1830_NOT));
and2 gate( .a(N3496_NOT), .b(p217), .O(EX541) );
and2 gate( .a(N1830_NOT), .b(EX541), .O(EX542) );
and2 gate( .a(N3496), .b(p218), .O(EX543) );
and2 gate( .a(N1830_NOT), .b(EX543), .O(EX544) );
and2 gate( .a(N3496_NOT), .b(p219), .O(EX545) );
and2 gate( .a(N1830), .b(EX545), .O(EX546) );
and2 gate( .a(N3496), .b(p220), .O(EX547) );
and2 gate( .a(N1830), .b(EX547), .O(EX548) );
or2  gate( .a(EX542), .b(EX544), .O(EX549) );
or2  gate( .a(EX546), .b(EX549), .O(EX550) );
or2  gate( .a(EX548), .b(EX550), .O(N4469) );
inv1 gate938( .a(N3496), .O(N4470) );
nand2 gate939( .a(N3499), .b(N1833), .O(N4471) );
inv1 gate940( .a(N3499), .O(N4472) );
inv1 gate941( .a(N3122), .O(N4473) );
inv1 gate942( .a(N3126), .O(N4474) );
nand2 gate943( .a(N3518), .b(N1840), .O(N4475) );
inv1 gate944( .a(N3518), .O(N4476) );
nand2 gate945( .a(N3521), .b(N1841), .O(N4477) );
inv1 gate946( .a(N3521), .O(N4478) );
nand2 gate947( .a(N3524), .b(N2275), .O(N4479) );
inv1 gate948( .a(N3524), .O(N4480) );
nand2 gate949( .a(N3527), .b(N1842), .O(N4481) );
inv1 gate950( .a(N3527), .O(N4482) );
inv1 gate( .a(N3530),.O(N3530_NOT) );
inv1 gate( .a(N1843),.O(N1843_NOT));
and2 gate( .a(N3530_NOT), .b(p221), .O(EX551) );
and2 gate( .a(N1843_NOT), .b(EX551), .O(EX552) );
and2 gate( .a(N3530), .b(p222), .O(EX553) );
and2 gate( .a(N1843_NOT), .b(EX553), .O(EX554) );
and2 gate( .a(N3530_NOT), .b(p223), .O(EX555) );
and2 gate( .a(N1843), .b(EX555), .O(EX556) );
and2 gate( .a(N3530), .b(p224), .O(EX557) );
and2 gate( .a(N1843), .b(EX557), .O(EX558) );
or2  gate( .a(EX552), .b(EX554), .O(EX559) );
or2  gate( .a(EX556), .b(EX559), .O(EX560) );
or2  gate( .a(EX558), .b(EX560), .O(N4483) );
inv1 gate952( .a(N3530), .O(N4484) );
inv1 gate953( .a(N3155), .O(N4485) );
inv1 gate954( .a(N3159), .O(N4486) );
nand2 gate955( .a(N1721), .b(N3954), .O(N4487) );
nand2 gate956( .a(N2235), .b(N3956), .O(N4488) );
inv1 gate957( .a(N3535), .O(N4489) );
nand2 gate958( .a(N3535), .b(N3958), .O(N4490) );
inv1 gate959( .a(N3539), .O(N4491) );
inv1 gate960( .a(N3542), .O(N4492) );
inv1 gate961( .a(N3545), .O(N4493) );
inv1 gate962( .a(N3548), .O(N4494) );
inv1 gate963( .a(N3553), .O(N4495) );
nand2 gate964( .a(N3553), .b(N3964), .O(N4496) );
inv1 gate965( .a(N3557), .O(N4497) );
inv1 gate966( .a(N3560), .O(N4498) );
inv1 gate967( .a(N3563), .O(N4499) );
inv1 gate968( .a(N3566), .O(N4500) );
inv1 gate969( .a(N3571), .O(N4501) );
nand2 gate970( .a(N3571), .b(N3167), .O(N4502) );
inv1 gate971( .a(N3574), .O(N4503) );
inv1 gate972( .a(N3577), .O(N4504) );
inv1 gate973( .a(N3580), .O(N4505) );
inv1 gate974( .a(N3583), .O(N4506) );
nand2 gate975( .a(N3598), .b(N1867), .O(N4507) );
inv1 gate976( .a(N3598), .O(N4508) );
nand2 gate977( .a(N3601), .b(N1868), .O(N4509) );
inv1 gate978( .a(N3601), .O(N4510) );
nand2 gate979( .a(N3604), .b(N1869), .O(N4511) );
inv1 gate980( .a(N3604), .O(N4512) );
nand2 gate981( .a(N3607), .b(N1870), .O(N4513) );
inv1 gate982( .a(N3607), .O(N4514) );
nand2 gate983( .a(N3610), .b(N1871), .O(N4515) );
inv1 gate984( .a(N3610), .O(N4516) );
nand2 gate985( .a(N3613), .b(N1872), .O(N4517) );
inv1 gate986( .a(N3613), .O(N4518) );
nand2 gate987( .a(N3616), .b(N1873), .O(N4519) );
inv1 gate988( .a(N3616), .O(N4520) );
nand2 gate989( .a(N3619), .b(N1874), .O(N4521) );
inv1 gate990( .a(N3619), .O(N4522) );
nand2 gate991( .a(N3622), .b(N1875), .O(N4523) );
inv1 gate992( .a(N3622), .O(N4524) );
nand2 gate993( .a(N3631), .b(N1876), .O(N4525) );
inv1 gate994( .a(N3631), .O(N4526) );
nand2 gate995( .a(N3634), .b(N1877), .O(N4527) );
inv1 gate996( .a(N3634), .O(N4528) );
nand2 gate997( .a(N3637), .b(N1878), .O(N4529) );
inv1 gate998( .a(N3637), .O(N4530) );
nand2 gate999( .a(N3640), .b(N1879), .O(N4531) );
inv1 gate1000( .a(N3640), .O(N4532) );
nand2 gate1001( .a(N3643), .b(N1880), .O(N4533) );
inv1 gate1002( .a(N3643), .O(N4534) );
nand2 gate1003( .a(N3646), .b(N1881), .O(N4535) );
inv1 gate1004( .a(N3646), .O(N4536) );
nand2 gate1005( .a(N3649), .b(N1882), .O(N4537) );
inv1 gate1006( .a(N3649), .O(N4538) );
inv1 gate( .a(N3652),.O(N3652_NOT) );
inv1 gate( .a(N1883),.O(N1883_NOT));
and2 gate( .a(N3652_NOT), .b(p225), .O(EX561) );
and2 gate( .a(N1883_NOT), .b(EX561), .O(EX562) );
and2 gate( .a(N3652), .b(p226), .O(EX563) );
and2 gate( .a(N1883_NOT), .b(EX563), .O(EX564) );
and2 gate( .a(N3652_NOT), .b(p227), .O(EX565) );
and2 gate( .a(N1883), .b(EX565), .O(EX566) );
and2 gate( .a(N3652), .b(p228), .O(EX567) );
and2 gate( .a(N1883), .b(EX567), .O(EX568) );
or2  gate( .a(EX562), .b(EX564), .O(EX569) );
or2  gate( .a(EX566), .b(EX569), .O(EX570) );
or2  gate( .a(EX568), .b(EX570), .O(N4539) );
inv1 gate1008( .a(N3652), .O(N4540) );
nand2 gate1009( .a(N3655), .b(N1884), .O(N4541) );
inv1 gate1010( .a(N3655), .O(N4542) );
inv1 gate1011( .a(N3658), .O(N4543) );
and2 gate1012( .a(N806), .b(N3293), .O(N4544) );
and2 gate1013( .a(N800), .b(N3287), .O(N4545) );
and2 gate1014( .a(N794), .b(N3281), .O(N4549) );
and2 gate1015( .a(N3273), .b(N786), .O(N4555) );
and2 gate1016( .a(N780), .b(N3267), .O(N4562) );
and2 gate1017( .a(N774), .b(N3355), .O(N4563) );
and2 gate1018( .a(N768), .b(N3349), .O(N4566) );
and2 gate1019( .a(N762), .b(N3343), .O(N4570) );
inv1 gate1020( .a(N3661), .O(N4575) );
inv1 gate( .a(N806),.O(N806_NOT) );
inv1 gate( .a(N3293),.O(N3293_NOT));
and2 gate( .a(N806_NOT), .b(p229), .O(EX571) );
and2 gate( .a(N3293_NOT), .b(EX571), .O(EX572) );
and2 gate( .a(N806), .b(p230), .O(EX573) );
and2 gate( .a(N3293_NOT), .b(EX573), .O(EX574) );
and2 gate( .a(N806_NOT), .b(p231), .O(EX575) );
and2 gate( .a(N3293), .b(EX575), .O(EX576) );
and2 gate( .a(N806), .b(p232), .O(EX577) );
and2 gate( .a(N3293), .b(EX577), .O(EX578) );
or2  gate( .a(EX572), .b(EX574), .O(EX579) );
or2  gate( .a(EX576), .b(EX579), .O(EX580) );
or2  gate( .a(EX578), .b(EX580), .O(N4576) );
and2 gate1022( .a(N800), .b(N3287), .O(N4577) );
and2 gate1023( .a(N794), .b(N3281), .O(N4581) );
and2 gate1024( .a(N786), .b(N3273), .O(N4586) );
and2 gate1025( .a(N780), .b(N3267), .O(N4592) );
and2 gate1026( .a(N774), .b(N3355), .O(N4593) );
and2 gate1027( .a(N768), .b(N3349), .O(N4597) );
and2 gate1028( .a(N762), .b(N3343), .O(N4603) );
inv1 gate1029( .a(N3664), .O(N4610) );
inv1 gate1030( .a(N3667), .O(N4611) );
inv1 gate1031( .a(N3670), .O(N4612) );
inv1 gate1032( .a(N3673), .O(N4613) );
inv1 gate1033( .a(N3676), .O(N4614) );
inv1 gate1034( .a(N3679), .O(N4615) );
inv1 gate1035( .a(N3682), .O(N4616) );
inv1 gate1036( .a(N3685), .O(N4617) );
inv1 gate1037( .a(N3688), .O(N4618) );
inv1 gate1038( .a(N3691), .O(N4619) );
inv1 gate1039( .a(N3694), .O(N4620) );
inv1 gate1040( .a(N3697), .O(N4621) );
inv1 gate1041( .a(N3700), .O(N4622) );
inv1 gate1042( .a(N3703), .O(N4623) );
inv1 gate1043( .a(N3706), .O(N4624) );
inv1 gate1044( .a(N3709), .O(N4625) );
inv1 gate1045( .a(N3712), .O(N4626) );
inv1 gate1046( .a(N3715), .O(N4627) );
inv1 gate1047( .a(N3718), .O(N4628) );
inv1 gate1048( .a(N3721), .O(N4629) );
and2 gate1049( .a(N3448), .b(N2704), .O(N4630) );
inv1 gate1050( .a(N3724), .O(N4631) );
and2 gate1051( .a(N3444), .b(N2700), .O(N4632) );
inv1 gate1052( .a(N3727), .O(N4633) );
and2 gate1053( .a(N3440), .b(N2696), .O(N4634) );
and2 gate1054( .a(N3436), .b(N2692), .O(N4635) );
inv1 gate1055( .a(N3730), .O(N4636) );
and2 gate1056( .a(N3432), .b(N2688), .O(N4637) );
and2 gate1057( .a(N3428), .b(N3311), .O(N4638) );
and2 gate1058( .a(N3424), .b(N3307), .O(N4639) );
and2 gate1059( .a(N3420), .b(N3303), .O(N4640) );
and2 gate1060( .a(N3416), .b(N3299), .O(N4641) );
inv1 gate1061( .a(N3733), .O(N4642) );
inv1 gate1062( .a(N3736), .O(N4643) );
inv1 gate1063( .a(N3739), .O(N4644) );
inv1 gate1064( .a(N3742), .O(N4645) );
inv1 gate1065( .a(N3745), .O(N4646) );
inv1 gate1066( .a(N3748), .O(N4647) );
inv1 gate1067( .a(N3751), .O(N4648) );
inv1 gate1068( .a(N3754), .O(N4649) );
inv1 gate1069( .a(N3757), .O(N4650) );
inv1 gate1070( .a(N3760), .O(N4651) );
inv1 gate1071( .a(N3763), .O(N4652) );
inv1 gate1072( .a(N3375), .O(N4653) );
and2 gate1073( .a(N865), .b(N3410), .O(N4656) );
inv1 gate( .a(N859),.O(N859_NOT) );
inv1 gate( .a(N3404),.O(N3404_NOT));
and2 gate( .a(N859_NOT), .b(p233), .O(EX581) );
and2 gate( .a(N3404_NOT), .b(EX581), .O(EX582) );
and2 gate( .a(N859), .b(p234), .O(EX583) );
and2 gate( .a(N3404_NOT), .b(EX583), .O(EX584) );
and2 gate( .a(N859_NOT), .b(p235), .O(EX585) );
and2 gate( .a(N3404), .b(EX585), .O(EX586) );
and2 gate( .a(N859), .b(p236), .O(EX587) );
and2 gate( .a(N3404), .b(EX587), .O(EX588) );
or2  gate( .a(EX582), .b(EX584), .O(EX589) );
or2  gate( .a(EX586), .b(EX589), .O(EX590) );
or2  gate( .a(EX588), .b(EX590), .O(N4657) );
and2 gate1075( .a(N853), .b(N3398), .O(N4661) );
and2 gate1076( .a(N3390), .b(N845), .O(N4667) );
and2 gate1077( .a(N839), .b(N3384), .O(N4674) );
and2 gate1078( .a(N833), .b(N3334), .O(N4675) );
and2 gate1079( .a(N827), .b(N3328), .O(N4678) );
and2 gate1080( .a(N821), .b(N3322), .O(N4682) );
and2 gate1081( .a(N814), .b(N3315), .O(N4687) );
inv1 gate1082( .a(N3766), .O(N4693) );
nand2 gate1083( .a(N3766), .b(N3380), .O(N4694) );
inv1 gate1084( .a(N3769), .O(N4695) );
inv1 gate1085( .a(N3772), .O(N4696) );
inv1 gate1086( .a(N3775), .O(N4697) );
inv1 gate1087( .a(N3778), .O(N4698) );
inv1 gate1088( .a(N3783), .O(N4699) );
inv1 gate1089( .a(N3786), .O(N4700) );
and2 gate1090( .a(N865), .b(N3410), .O(N4701) );
and2 gate1091( .a(N859), .b(N3404), .O(N4702) );
and2 gate1092( .a(N853), .b(N3398), .O(N4706) );
and2 gate1093( .a(N845), .b(N3390), .O(N4711) );
and2 gate1094( .a(N839), .b(N3384), .O(N4717) );
and2 gate1095( .a(N833), .b(N3334), .O(N4718) );
and2 gate1096( .a(N827), .b(N3328), .O(N4722) );
and2 gate1097( .a(N821), .b(N3322), .O(N4728) );
and2 gate1098( .a(N814), .b(N3315), .O(N4735) );
inv1 gate1099( .a(N3789), .O(N4743) );
inv1 gate1100( .a(N3792), .O(N4744) );
inv1 gate1101( .a(N3807), .O(N4745) );
nand2 gate1102( .a(N3807), .b(N3452), .O(N4746) );
inv1 gate1103( .a(N3810), .O(N4747) );
inv1 gate1104( .a(N3813), .O(N4748) );
inv1 gate1105( .a(N3816), .O(N4749) );
inv1 gate1106( .a(N3819), .O(N4750) );
nand2 gate1107( .a(N3819), .b(N3453), .O(N4751) );
inv1 gate1108( .a(N3822), .O(N4752) );
inv1 gate1109( .a(N3825), .O(N4753) );
inv1 gate1110( .a(N3828), .O(N4754) );
inv1 gate1111( .a(N3831), .O(N4755) );
and2 gate1112( .a(N3482), .b(N3263), .O(N4756) );
and2 gate1113( .a(N3478), .b(N3259), .O(N4757) );
and2 gate1114( .a(N3474), .b(N3255), .O(N4758) );
and2 gate1115( .a(N3470), .b(N3251), .O(N4759) );
and2 gate1116( .a(N3466), .b(N3247), .O(N4760) );
inv1 gate1117( .a(N3846), .O(N4761) );
and2 gate1118( .a(N3462), .b(N2615), .O(N4762) );
inv1 gate1119( .a(N3849), .O(N4763) );
and2 gate1120( .a(N3458), .b(N2611), .O(N4764) );
inv1 gate1121( .a(N3852), .O(N4765) );
and2 gate1122( .a(N3454), .b(N2607), .O(N4766) );
and2 gate1123( .a(N2680), .b(N3381), .O(N4767) );
inv1 gate1124( .a(N3855), .O(N4768) );
and2 gate1125( .a(N3340), .b(N695), .O(N4769) );
inv1 gate1126( .a(N3858), .O(N4775) );
inv1 gate( .a(N3858),.O(N3858_NOT) );
inv1 gate( .a(N3486),.O(N3486_NOT));
and2 gate( .a(N3858_NOT), .b(p237), .O(EX591) );
and2 gate( .a(N3486_NOT), .b(EX591), .O(EX592) );
and2 gate( .a(N3858), .b(p238), .O(EX593) );
and2 gate( .a(N3486_NOT), .b(EX593), .O(EX594) );
and2 gate( .a(N3858_NOT), .b(p239), .O(EX595) );
and2 gate( .a(N3486), .b(EX595), .O(EX596) );
and2 gate( .a(N3858), .b(p240), .O(EX597) );
and2 gate( .a(N3486), .b(EX597), .O(EX598) );
or2  gate( .a(EX592), .b(EX594), .O(EX599) );
or2  gate( .a(EX596), .b(EX599), .O(EX600) );
or2  gate( .a(EX598), .b(EX600), .O(N4776) );
inv1 gate1128( .a(N3861), .O(N4777) );
inv1 gate1129( .a(N3864), .O(N4778) );
inv1 gate1130( .a(N3867), .O(N4779) );
inv1 gate1131( .a(N3870), .O(N4780) );
inv1 gate1132( .a(N3885), .O(N4781) );
inv1 gate1133( .a(N3888), .O(N4782) );
inv1 gate1134( .a(N3891), .O(N4783) );
or2 gate1135( .a(N3131), .b(N3134), .O(N4784) );
inv1 gate1136( .a(N3502), .O(N4789) );
inv1 gate1137( .a(N3131), .O(N4790) );
inv1 gate1138( .a(N3507), .O(N4793) );
inv1 gate1139( .a(N3510), .O(N4794) );
inv1 gate1140( .a(N3515), .O(N4795) );
buf1 gate1141( .a(N3114), .O(N4796) );
inv1 gate1142( .a(N3586), .O(N4799) );
inv1 gate1143( .a(N3589), .O(N4800) );
inv1 gate1144( .a(N3592), .O(N4801) );
inv1 gate1145( .a(N3595), .O(N4802) );
nand2 gate1146( .a(N4326), .b(N4327), .O(N4803) );
inv1 gate( .a(N4333),.O(N4333_NOT) );
inv1 gate( .a(N4334),.O(N4334_NOT));
and2 gate( .a(N4333_NOT), .b(p241), .O(EX601) );
and2 gate( .a(N4334_NOT), .b(EX601), .O(EX602) );
and2 gate( .a(N4333), .b(p242), .O(EX603) );
and2 gate( .a(N4334_NOT), .b(EX603), .O(EX604) );
and2 gate( .a(N4333_NOT), .b(p243), .O(EX605) );
and2 gate( .a(N4334), .b(EX605), .O(EX606) );
and2 gate( .a(N4333), .b(p244), .O(EX607) );
and2 gate( .a(N4334), .b(EX607), .O(EX608) );
or2  gate( .a(EX602), .b(EX604), .O(EX609) );
or2  gate( .a(EX606), .b(EX609), .O(EX610) );
or2  gate( .a(EX608), .b(EX610), .O(N4806) );
inv1 gate1148( .a(N3625), .O(N4809) );
buf1 gate1149( .a(N3178), .O(N4810) );
inv1 gate1150( .a(N3628), .O(N4813) );
buf1 gate1151( .a(N3202), .O(N4814) );
buf1 gate1152( .a(N3221), .O(N4817) );
buf1 gate1153( .a(N3293), .O(N4820) );
buf1 gate1154( .a(N3287), .O(N4823) );
buf1 gate1155( .a(N3281), .O(N4826) );
buf1 gate1156( .a(N3273), .O(N4829) );
buf1 gate1157( .a(N3267), .O(N4832) );
buf1 gate1158( .a(N3355), .O(N4835) );
buf1 gate1159( .a(N3349), .O(N4838) );
buf1 gate1160( .a(N3343), .O(N4841) );
nor2 gate1161( .a(N3273), .b(N786), .O(N4844) );
buf1 gate1162( .a(N3293), .O(N4847) );
buf1 gate1163( .a(N3287), .O(N4850) );
buf1 gate1164( .a(N3281), .O(N4853) );
buf1 gate1165( .a(N3267), .O(N4856) );
buf1 gate1166( .a(N3355), .O(N4859) );
buf1 gate1167( .a(N3349), .O(N4862) );
buf1 gate1168( .a(N3343), .O(N4865) );
buf1 gate1169( .a(N3273), .O(N4868) );
nor2 gate1170( .a(N786), .b(N3273), .O(N4871) );
buf1 gate1171( .a(N3448), .O(N4874) );
buf1 gate1172( .a(N3444), .O(N4877) );
buf1 gate1173( .a(N3440), .O(N4880) );
buf1 gate1174( .a(N3432), .O(N4883) );
buf1 gate1175( .a(N3428), .O(N4886) );
buf1 gate1176( .a(N3311), .O(N4889) );
buf1 gate1177( .a(N3424), .O(N4892) );
buf1 gate1178( .a(N3307), .O(N4895) );
buf1 gate1179( .a(N3420), .O(N4898) );
buf1 gate1180( .a(N3303), .O(N4901) );
buf1 gate1181( .a(N3436), .O(N4904) );
buf1 gate1182( .a(N3416), .O(N4907) );
buf1 gate1183( .a(N3299), .O(N4910) );
buf1 gate1184( .a(N3410), .O(N4913) );
buf1 gate1185( .a(N3404), .O(N4916) );
buf1 gate1186( .a(N3398), .O(N4919) );
buf1 gate1187( .a(N3390), .O(N4922) );
buf1 gate1188( .a(N3384), .O(N4925) );
buf1 gate1189( .a(N3334), .O(N4928) );
buf1 gate1190( .a(N3328), .O(N4931) );
buf1 gate1191( .a(N3322), .O(N4934) );
buf1 gate1192( .a(N3315), .O(N4937) );
nor2 gate1193( .a(N3390), .b(N845), .O(N4940) );
buf1 gate1194( .a(N3315), .O(N4943) );
buf1 gate1195( .a(N3328), .O(N4946) );
buf1 gate1196( .a(N3322), .O(N4949) );
buf1 gate1197( .a(N3384), .O(N4952) );
buf1 gate1198( .a(N3334), .O(N4955) );
buf1 gate1199( .a(N3398), .O(N4958) );
buf1 gate1200( .a(N3390), .O(N4961) );
buf1 gate1201( .a(N3410), .O(N4964) );
buf1 gate1202( .a(N3404), .O(N4967) );
buf1 gate1203( .a(N3340), .O(N4970) );
buf1 gate1204( .a(N3349), .O(N4973) );
buf1 gate1205( .a(N3343), .O(N4976) );
buf1 gate1206( .a(N3267), .O(N4979) );
buf1 gate1207( .a(N3355), .O(N4982) );
buf1 gate1208( .a(N3281), .O(N4985) );
buf1 gate1209( .a(N3273), .O(N4988) );
buf1 gate1210( .a(N3293), .O(N4991) );
buf1 gate1211( .a(N3287), .O(N4994) );
nand2 gate1212( .a(N4411), .b(N4412), .O(N4997) );
buf1 gate1213( .a(N3410), .O(N5000) );
buf1 gate1214( .a(N3404), .O(N5003) );
buf1 gate1215( .a(N3398), .O(N5006) );
buf1 gate1216( .a(N3384), .O(N5009) );
buf1 gate1217( .a(N3334), .O(N5012) );
buf1 gate1218( .a(N3328), .O(N5015) );
buf1 gate1219( .a(N3322), .O(N5018) );
buf1 gate1220( .a(N3390), .O(N5021) );
buf1 gate1221( .a(N3315), .O(N5024) );
nor2 gate1222( .a(N845), .b(N3390), .O(N5027) );
nor2 gate1223( .a(N814), .b(N3315), .O(N5030) );
buf1 gate1224( .a(N3299), .O(N5033) );
buf1 gate1225( .a(N3307), .O(N5036) );
buf1 gate1226( .a(N3303), .O(N5039) );
buf1 gate1227( .a(N3311), .O(N5042) );
inv1 gate1228( .a(N3795), .O(N5045) );
inv1 gate1229( .a(N3798), .O(N5046) );
inv1 gate1230( .a(N3801), .O(N5047) );
inv1 gate1231( .a(N3804), .O(N5048) );
buf1 gate1232( .a(N3247), .O(N5049) );
buf1 gate1233( .a(N3255), .O(N5052) );
buf1 gate1234( .a(N3251), .O(N5055) );
buf1 gate1235( .a(N3263), .O(N5058) );
buf1 gate1236( .a(N3259), .O(N5061) );
inv1 gate1237( .a(N3834), .O(N5064) );
inv1 gate1238( .a(N3837), .O(N5065) );
inv1 gate1239( .a(N3840), .O(N5066) );
inv1 gate1240( .a(N3843), .O(N5067) );
buf1 gate1241( .a(N3482), .O(N5068) );
buf1 gate1242( .a(N3263), .O(N5071) );
buf1 gate1243( .a(N3478), .O(N5074) );
buf1 gate1244( .a(N3259), .O(N5077) );
buf1 gate1245( .a(N3474), .O(N5080) );
buf1 gate1246( .a(N3255), .O(N5083) );
buf1 gate1247( .a(N3466), .O(N5086) );
buf1 gate1248( .a(N3247), .O(N5089) );
buf1 gate1249( .a(N3462), .O(N5092) );
buf1 gate1250( .a(N3458), .O(N5095) );
buf1 gate1251( .a(N3454), .O(N5098) );
buf1 gate1252( .a(N3470), .O(N5101) );
buf1 gate1253( .a(N3251), .O(N5104) );
buf1 gate1254( .a(N3381), .O(N5107) );
inv1 gate1255( .a(N3873), .O(N5110) );
inv1 gate1256( .a(N3876), .O(N5111) );
inv1 gate1257( .a(N3879), .O(N5112) );
inv1 gate1258( .a(N3882), .O(N5113) );
buf1 gate1259( .a(N3458), .O(N5114) );
buf1 gate1260( .a(N3454), .O(N5117) );
buf1 gate1261( .a(N3466), .O(N5120) );
buf1 gate1262( .a(N3462), .O(N5123) );
buf1 gate1263( .a(N3474), .O(N5126) );
buf1 gate1264( .a(N3470), .O(N5129) );
buf1 gate1265( .a(N3482), .O(N5132) );
buf1 gate1266( .a(N3478), .O(N5135) );
buf1 gate1267( .a(N3416), .O(N5138) );
buf1 gate1268( .a(N3424), .O(N5141) );
buf1 gate1269( .a(N3420), .O(N5144) );
buf1 gate1270( .a(N3432), .O(N5147) );
buf1 gate1271( .a(N3428), .O(N5150) );
buf1 gate1272( .a(N3440), .O(N5153) );
buf1 gate1273( .a(N3436), .O(N5156) );
buf1 gate1274( .a(N3448), .O(N5159) );
buf1 gate1275( .a(N3444), .O(N5162) );
nand2 gate1276( .a(N4486), .b(N4485), .O(N5165) );
nand2 gate1277( .a(N4474), .b(N4473), .O(N5166) );
nand2 gate1278( .a(N1290), .b(N4464), .O(N5167) );
nand2 gate1279( .a(N1293), .b(N4466), .O(N5168) );
nand2 gate1280( .a(N2074), .b(N4468), .O(N5169) );
nand2 gate1281( .a(N1296), .b(N4470), .O(N5170) );
nand2 gate1282( .a(N1302), .b(N4472), .O(N5171) );
nand2 gate1283( .a(N1314), .b(N4476), .O(N5172) );
nand2 gate1284( .a(N1317), .b(N4478), .O(N5173) );
nand2 gate1285( .a(N2081), .b(N4480), .O(N5174) );
nand2 gate1286( .a(N1320), .b(N4482), .O(N5175) );
nand2 gate1287( .a(N1323), .b(N4484), .O(N5176) );
nand2 gate1288( .a(N3953), .b(N4487), .O(N5177) );
nand2 gate1289( .a(N3955), .b(N4488), .O(N5178) );
nand2 gate1290( .a(N3073), .b(N4489), .O(N5179) );
nand2 gate1291( .a(N3542), .b(N4491), .O(N5180) );
nand2 gate1292( .a(N3539), .b(N4492), .O(N5181) );
nand2 gate1293( .a(N3548), .b(N4493), .O(N5182) );
inv1 gate( .a(N3545),.O(N3545_NOT) );
inv1 gate( .a(N4494),.O(N4494_NOT));
and2 gate( .a(N3545_NOT), .b(p245), .O(EX611) );
and2 gate( .a(N4494_NOT), .b(EX611), .O(EX612) );
and2 gate( .a(N3545), .b(p246), .O(EX613) );
and2 gate( .a(N4494_NOT), .b(EX613), .O(EX614) );
and2 gate( .a(N3545_NOT), .b(p247), .O(EX615) );
and2 gate( .a(N4494), .b(EX615), .O(EX616) );
and2 gate( .a(N3545), .b(p248), .O(EX617) );
and2 gate( .a(N4494), .b(EX617), .O(EX618) );
or2  gate( .a(EX612), .b(EX614), .O(EX619) );
or2  gate( .a(EX616), .b(EX619), .O(EX620) );
or2  gate( .a(EX618), .b(EX620), .O(N5183) );
nand2 gate1295( .a(N3080), .b(N4495), .O(N5184) );
nand2 gate1296( .a(N3560), .b(N4497), .O(N5185) );
nand2 gate1297( .a(N3557), .b(N4498), .O(N5186) );
nand2 gate1298( .a(N3566), .b(N4499), .O(N5187) );
inv1 gate( .a(N3563),.O(N3563_NOT) );
inv1 gate( .a(N4500),.O(N4500_NOT));
and2 gate( .a(N3563_NOT), .b(p249), .O(EX621) );
and2 gate( .a(N4500_NOT), .b(EX621), .O(EX622) );
and2 gate( .a(N3563), .b(p250), .O(EX623) );
and2 gate( .a(N4500_NOT), .b(EX623), .O(EX624) );
and2 gate( .a(N3563_NOT), .b(p251), .O(EX625) );
and2 gate( .a(N4500), .b(EX625), .O(EX626) );
and2 gate( .a(N3563), .b(p252), .O(EX627) );
and2 gate( .a(N4500), .b(EX627), .O(EX628) );
or2  gate( .a(EX622), .b(EX624), .O(EX629) );
or2  gate( .a(EX626), .b(EX629), .O(EX630) );
or2  gate( .a(EX628), .b(EX630), .O(N5188) );
nand2 gate1300( .a(N2778), .b(N4501), .O(N5189) );
nand2 gate1301( .a(N3577), .b(N4503), .O(N5190) );
nand2 gate1302( .a(N3574), .b(N4504), .O(N5191) );
nand2 gate1303( .a(N3583), .b(N4505), .O(N5192) );
nand2 gate1304( .a(N3580), .b(N4506), .O(N5193) );
nand2 gate1305( .a(N1326), .b(N4508), .O(N5196) );
nand2 gate1306( .a(N1329), .b(N4510), .O(N5197) );
nand2 gate1307( .a(N1332), .b(N4512), .O(N5198) );
nand2 gate1308( .a(N1335), .b(N4514), .O(N5199) );
nand2 gate1309( .a(N1338), .b(N4516), .O(N5200) );
nand2 gate1310( .a(N1341), .b(N4518), .O(N5201) );
nand2 gate1311( .a(N1344), .b(N4520), .O(N5202) );
nand2 gate1312( .a(N1347), .b(N4522), .O(N5203) );
nand2 gate1313( .a(N1350), .b(N4524), .O(N5204) );
nand2 gate1314( .a(N1353), .b(N4526), .O(N5205) );
nand2 gate1315( .a(N1356), .b(N4528), .O(N5206) );
nand2 gate1316( .a(N1359), .b(N4530), .O(N5207) );
nand2 gate1317( .a(N1362), .b(N4532), .O(N5208) );
nand2 gate1318( .a(N1365), .b(N4534), .O(N5209) );
inv1 gate( .a(N1368),.O(N1368_NOT) );
inv1 gate( .a(N4536),.O(N4536_NOT));
and2 gate( .a(N1368_NOT), .b(p253), .O(EX631) );
and2 gate( .a(N4536_NOT), .b(EX631), .O(EX632) );
and2 gate( .a(N1368), .b(p254), .O(EX633) );
and2 gate( .a(N4536_NOT), .b(EX633), .O(EX634) );
and2 gate( .a(N1368_NOT), .b(p255), .O(EX635) );
and2 gate( .a(N4536), .b(EX635), .O(EX636) );
and2 gate( .a(N1368), .b(p256), .O(EX637) );
and2 gate( .a(N4536), .b(EX637), .O(EX638) );
or2  gate( .a(EX632), .b(EX634), .O(EX639) );
or2  gate( .a(EX636), .b(EX639), .O(EX640) );
or2  gate( .a(EX638), .b(EX640), .O(N5210) );
nand2 gate1320( .a(N1371), .b(N4538), .O(N5211) );
nand2 gate1321( .a(N1374), .b(N4540), .O(N5212) );
nand2 gate1322( .a(N1377), .b(N4542), .O(N5213) );
inv1 gate( .a(N3670),.O(N3670_NOT) );
inv1 gate( .a(N4611),.O(N4611_NOT));
and2 gate( .a(N3670_NOT), .b(p257), .O(EX641) );
and2 gate( .a(N4611_NOT), .b(EX641), .O(EX642) );
and2 gate( .a(N3670), .b(p258), .O(EX643) );
and2 gate( .a(N4611_NOT), .b(EX643), .O(EX644) );
and2 gate( .a(N3670_NOT), .b(p259), .O(EX645) );
and2 gate( .a(N4611), .b(EX645), .O(EX646) );
and2 gate( .a(N3670), .b(p260), .O(EX647) );
and2 gate( .a(N4611), .b(EX647), .O(EX648) );
or2  gate( .a(EX642), .b(EX644), .O(EX649) );
or2  gate( .a(EX646), .b(EX649), .O(EX650) );
or2  gate( .a(EX648), .b(EX650), .O(N5283) );
nand2 gate1324( .a(N3667), .b(N4612), .O(N5284) );
nand2 gate1325( .a(N3676), .b(N4613), .O(N5285) );
nand2 gate1326( .a(N3673), .b(N4614), .O(N5286) );
nand2 gate1327( .a(N3682), .b(N4615), .O(N5287) );
nand2 gate1328( .a(N3679), .b(N4616), .O(N5288) );
nand2 gate1329( .a(N3688), .b(N4617), .O(N5289) );
nand2 gate1330( .a(N3685), .b(N4618), .O(N5290) );
nand2 gate1331( .a(N3694), .b(N4619), .O(N5291) );
nand2 gate1332( .a(N3691), .b(N4620), .O(N5292) );
nand2 gate1333( .a(N3700), .b(N4621), .O(N5293) );
nand2 gate1334( .a(N3697), .b(N4622), .O(N5294) );
nand2 gate1335( .a(N3706), .b(N4623), .O(N5295) );
nand2 gate1336( .a(N3703), .b(N4624), .O(N5296) );
nand2 gate1337( .a(N3712), .b(N4625), .O(N5297) );
nand2 gate1338( .a(N3709), .b(N4626), .O(N5298) );
nand2 gate1339( .a(N3718), .b(N4627), .O(N5299) );
nand2 gate1340( .a(N3715), .b(N4628), .O(N5300) );
nand2 gate1341( .a(N3739), .b(N4643), .O(N5314) );
nand2 gate1342( .a(N3736), .b(N4644), .O(N5315) );
nand2 gate1343( .a(N3745), .b(N4645), .O(N5316) );
nand2 gate1344( .a(N3742), .b(N4646), .O(N5317) );
inv1 gate( .a(N3751),.O(N3751_NOT) );
inv1 gate( .a(N4647),.O(N4647_NOT));
and2 gate( .a(N3751_NOT), .b(p261), .O(EX651) );
and2 gate( .a(N4647_NOT), .b(EX651), .O(EX652) );
and2 gate( .a(N3751), .b(p262), .O(EX653) );
and2 gate( .a(N4647_NOT), .b(EX653), .O(EX654) );
and2 gate( .a(N3751_NOT), .b(p263), .O(EX655) );
and2 gate( .a(N4647), .b(EX655), .O(EX656) );
and2 gate( .a(N3751), .b(p264), .O(EX657) );
and2 gate( .a(N4647), .b(EX657), .O(EX658) );
or2  gate( .a(EX652), .b(EX654), .O(EX659) );
or2  gate( .a(EX656), .b(EX659), .O(EX660) );
or2  gate( .a(EX658), .b(EX660), .O(N5318) );
nand2 gate1346( .a(N3748), .b(N4648), .O(N5319) );
nand2 gate1347( .a(N3757), .b(N4649), .O(N5320) );
inv1 gate( .a(N3754),.O(N3754_NOT) );
inv1 gate( .a(N4650),.O(N4650_NOT));
and2 gate( .a(N3754_NOT), .b(p265), .O(EX661) );
and2 gate( .a(N4650_NOT), .b(EX661), .O(EX662) );
and2 gate( .a(N3754), .b(p266), .O(EX663) );
and2 gate( .a(N4650_NOT), .b(EX663), .O(EX664) );
and2 gate( .a(N3754_NOT), .b(p267), .O(EX665) );
and2 gate( .a(N4650), .b(EX665), .O(EX666) );
and2 gate( .a(N3754), .b(p268), .O(EX667) );
and2 gate( .a(N4650), .b(EX667), .O(EX668) );
or2  gate( .a(EX662), .b(EX664), .O(EX669) );
or2  gate( .a(EX666), .b(EX669), .O(EX670) );
or2  gate( .a(EX668), .b(EX670), .O(N5321) );
nand2 gate1349( .a(N3763), .b(N4651), .O(N5322) );
inv1 gate( .a(N3760),.O(N3760_NOT) );
inv1 gate( .a(N4652),.O(N4652_NOT));
and2 gate( .a(N3760_NOT), .b(p269), .O(EX671) );
and2 gate( .a(N4652_NOT), .b(EX671), .O(EX672) );
and2 gate( .a(N3760), .b(p270), .O(EX673) );
and2 gate( .a(N4652_NOT), .b(EX673), .O(EX674) );
and2 gate( .a(N3760_NOT), .b(p271), .O(EX675) );
and2 gate( .a(N4652), .b(EX675), .O(EX676) );
and2 gate( .a(N3760), .b(p272), .O(EX677) );
and2 gate( .a(N4652), .b(EX677), .O(EX678) );
or2  gate( .a(EX672), .b(EX674), .O(EX679) );
or2  gate( .a(EX676), .b(EX679), .O(EX680) );
or2  gate( .a(EX678), .b(EX680), .O(N5323) );
inv1 gate1351( .a(N4193), .O(N5324) );
nand2 gate1352( .a(N2781), .b(N4693), .O(N5363) );
inv1 gate( .a(N3772),.O(N3772_NOT) );
inv1 gate( .a(N4695),.O(N4695_NOT));
and2 gate( .a(N3772_NOT), .b(p273), .O(EX681) );
and2 gate( .a(N4695_NOT), .b(EX681), .O(EX682) );
and2 gate( .a(N3772), .b(p274), .O(EX683) );
and2 gate( .a(N4695_NOT), .b(EX683), .O(EX684) );
and2 gate( .a(N3772_NOT), .b(p275), .O(EX685) );
and2 gate( .a(N4695), .b(EX685), .O(EX686) );
and2 gate( .a(N3772), .b(p276), .O(EX687) );
and2 gate( .a(N4695), .b(EX687), .O(EX688) );
or2  gate( .a(EX682), .b(EX684), .O(EX689) );
or2  gate( .a(EX686), .b(EX689), .O(EX690) );
or2  gate( .a(EX688), .b(EX690), .O(N5364) );
nand2 gate1354( .a(N3769), .b(N4696), .O(N5365) );
nand2 gate1355( .a(N3778), .b(N4697), .O(N5366) );
nand2 gate1356( .a(N3775), .b(N4698), .O(N5367) );
nand2 gate1357( .a(N2790), .b(N4745), .O(N5425) );
nand2 gate1358( .a(N3813), .b(N4747), .O(N5426) );
nand2 gate1359( .a(N3810), .b(N4748), .O(N5427) );
nand2 gate1360( .a(N2793), .b(N4750), .O(N5429) );
nand2 gate1361( .a(N3825), .b(N4752), .O(N5430) );
nand2 gate1362( .a(N3822), .b(N4753), .O(N5431) );
nand2 gate1363( .a(N3831), .b(N4754), .O(N5432) );
nand2 gate1364( .a(N3828), .b(N4755), .O(N5433) );
nand2 gate1365( .a(N2796), .b(N4775), .O(N5451) );
nand2 gate1366( .a(N3864), .b(N4777), .O(N5452) );
nand2 gate1367( .a(N3861), .b(N4778), .O(N5453) );
nand2 gate1368( .a(N3870), .b(N4779), .O(N5454) );
nand2 gate1369( .a(N3867), .b(N4780), .O(N5455) );
nand2 gate1370( .a(N3888), .b(N4781), .O(N5456) );
nand2 gate1371( .a(N3885), .b(N4782), .O(N5457) );
inv1 gate1372( .a(N4303), .O(N5469) );
nand2 gate1373( .a(N3589), .b(N4799), .O(N5474) );
nand2 gate1374( .a(N3586), .b(N4800), .O(N5475) );
nand2 gate1375( .a(N3595), .b(N4801), .O(N5476) );
nand2 gate1376( .a(N3592), .b(N4802), .O(N5477) );
inv1 gate( .a(N3798),.O(N3798_NOT) );
inv1 gate( .a(N5045),.O(N5045_NOT));
and2 gate( .a(N3798_NOT), .b(p277), .O(EX691) );
and2 gate( .a(N5045_NOT), .b(EX691), .O(EX692) );
and2 gate( .a(N3798), .b(p278), .O(EX693) );
and2 gate( .a(N5045_NOT), .b(EX693), .O(EX694) );
and2 gate( .a(N3798_NOT), .b(p279), .O(EX695) );
and2 gate( .a(N5045), .b(EX695), .O(EX696) );
and2 gate( .a(N3798), .b(p280), .O(EX697) );
and2 gate( .a(N5045), .b(EX697), .O(EX698) );
or2  gate( .a(EX692), .b(EX694), .O(EX699) );
or2  gate( .a(EX696), .b(EX699), .O(EX700) );
or2  gate( .a(EX698), .b(EX700), .O(N5571) );
nand2 gate1378( .a(N3795), .b(N5046), .O(N5572) );
nand2 gate1379( .a(N3804), .b(N5047), .O(N5573) );
nand2 gate1380( .a(N3801), .b(N5048), .O(N5574) );
nand2 gate1381( .a(N3837), .b(N5064), .O(N5584) );
nand2 gate1382( .a(N3834), .b(N5065), .O(N5585) );
nand2 gate1383( .a(N3843), .b(N5066), .O(N5586) );
nand2 gate1384( .a(N3840), .b(N5067), .O(N5587) );
nand2 gate1385( .a(N3876), .b(N5110), .O(N5602) );
nand2 gate1386( .a(N3873), .b(N5111), .O(N5603) );
nand2 gate1387( .a(N3882), .b(N5112), .O(N5604) );
nand2 gate1388( .a(N3879), .b(N5113), .O(N5605) );
nand2 gate1389( .a(N5324), .b(N4653), .O(N5631) );
nand2 gate1390( .a(N4463), .b(N5167), .O(N5632) );
nand2 gate1391( .a(N4465), .b(N5168), .O(N5640) );
nand2 gate1392( .a(N4467), .b(N5169), .O(N5654) );
nand2 gate1393( .a(N4469), .b(N5170), .O(N5670) );
nand2 gate1394( .a(N4471), .b(N5171), .O(N5683) );
nand2 gate1395( .a(N4475), .b(N5172), .O(N5690) );
nand2 gate1396( .a(N4477), .b(N5173), .O(N5697) );
nand2 gate1397( .a(N4479), .b(N5174), .O(N5707) );
inv1 gate( .a(N4481),.O(N4481_NOT) );
inv1 gate( .a(N5175),.O(N5175_NOT));
and2 gate( .a(N4481_NOT), .b(p281), .O(EX701) );
and2 gate( .a(N5175_NOT), .b(EX701), .O(EX702) );
and2 gate( .a(N4481), .b(p282), .O(EX703) );
and2 gate( .a(N5175_NOT), .b(EX703), .O(EX704) );
and2 gate( .a(N4481_NOT), .b(p283), .O(EX705) );
and2 gate( .a(N5175), .b(EX705), .O(EX706) );
and2 gate( .a(N4481), .b(p284), .O(EX707) );
and2 gate( .a(N5175), .b(EX707), .O(EX708) );
or2  gate( .a(EX702), .b(EX704), .O(EX709) );
or2  gate( .a(EX706), .b(EX709), .O(EX710) );
or2  gate( .a(EX708), .b(EX710), .O(N5718) );
nand2 gate1399( .a(N4483), .b(N5176), .O(N5728) );
inv1 gate1400( .a(N5177), .O(N5735) );
nand2 gate1401( .a(N5179), .b(N4490), .O(N5736) );
nand2 gate1402( .a(N5180), .b(N5181), .O(N5740) );
nand2 gate1403( .a(N5182), .b(N5183), .O(N5744) );
nand2 gate1404( .a(N5184), .b(N4496), .O(N5747) );
nand2 gate1405( .a(N5185), .b(N5186), .O(N5751) );
nand2 gate1406( .a(N5187), .b(N5188), .O(N5755) );
nand2 gate1407( .a(N5189), .b(N4502), .O(N5758) );
nand2 gate1408( .a(N5190), .b(N5191), .O(N5762) );
inv1 gate( .a(N5192),.O(N5192_NOT) );
inv1 gate( .a(N5193),.O(N5193_NOT));
and2 gate( .a(N5192_NOT), .b(p285), .O(EX711) );
and2 gate( .a(N5193_NOT), .b(EX711), .O(EX712) );
and2 gate( .a(N5192), .b(p286), .O(EX713) );
and2 gate( .a(N5193_NOT), .b(EX713), .O(EX714) );
and2 gate( .a(N5192_NOT), .b(p287), .O(EX715) );
and2 gate( .a(N5193), .b(EX715), .O(EX716) );
and2 gate( .a(N5192), .b(p288), .O(EX717) );
and2 gate( .a(N5193), .b(EX717), .O(EX718) );
or2  gate( .a(EX712), .b(EX714), .O(EX719) );
or2  gate( .a(EX716), .b(EX719), .O(EX720) );
or2  gate( .a(EX718), .b(EX720), .O(N5766) );
inv1 gate1410( .a(N4803), .O(N5769) );
inv1 gate1411( .a(N4806), .O(N5770) );
nand2 gate1412( .a(N4507), .b(N5196), .O(N5771) );
nand2 gate1413( .a(N4509), .b(N5197), .O(N5778) );
nand2 gate1414( .a(N4511), .b(N5198), .O(N5789) );
nand2 gate1415( .a(N4513), .b(N5199), .O(N5799) );
nand2 gate1416( .a(N4515), .b(N5200), .O(N5807) );
nand2 gate1417( .a(N4517), .b(N5201), .O(N5821) );
nand2 gate1418( .a(N4519), .b(N5202), .O(N5837) );
nand2 gate1419( .a(N4521), .b(N5203), .O(N5850) );
nand2 gate1420( .a(N4523), .b(N5204), .O(N5856) );
nand2 gate1421( .a(N4525), .b(N5205), .O(N5863) );
nand2 gate1422( .a(N4527), .b(N5206), .O(N5870) );
nand2 gate1423( .a(N4529), .b(N5207), .O(N5881) );
nand2 gate1424( .a(N4531), .b(N5208), .O(N5892) );
nand2 gate1425( .a(N4533), .b(N5209), .O(N5898) );
nand2 gate1426( .a(N4535), .b(N5210), .O(N5905) );
nand2 gate1427( .a(N4537), .b(N5211), .O(N5915) );
inv1 gate( .a(N4539),.O(N4539_NOT) );
inv1 gate( .a(N5212),.O(N5212_NOT));
and2 gate( .a(N4539_NOT), .b(p289), .O(EX721) );
and2 gate( .a(N5212_NOT), .b(EX721), .O(EX722) );
and2 gate( .a(N4539), .b(p290), .O(EX723) );
and2 gate( .a(N5212_NOT), .b(EX723), .O(EX724) );
and2 gate( .a(N4539_NOT), .b(p291), .O(EX725) );
and2 gate( .a(N5212), .b(EX725), .O(EX726) );
and2 gate( .a(N4539), .b(p292), .O(EX727) );
and2 gate( .a(N5212), .b(EX727), .O(EX728) );
or2  gate( .a(EX722), .b(EX724), .O(EX729) );
or2  gate( .a(EX726), .b(EX729), .O(EX730) );
or2  gate( .a(EX728), .b(EX730), .O(N5926) );
nand2 gate1429( .a(N4541), .b(N5213), .O(N5936) );
inv1 gate1430( .a(N4817), .O(N5943) );
nand2 gate1431( .a(N4820), .b(N1931), .O(N5944) );
inv1 gate1432( .a(N4820), .O(N5945) );
nand2 gate1433( .a(N4823), .b(N1932), .O(N5946) );
inv1 gate1434( .a(N4823), .O(N5947) );
nand2 gate1435( .a(N4826), .b(N1933), .O(N5948) );
inv1 gate1436( .a(N4826), .O(N5949) );
nand2 gate1437( .a(N4829), .b(N1934), .O(N5950) );
inv1 gate1438( .a(N4829), .O(N5951) );
nand2 gate1439( .a(N4832), .b(N1935), .O(N5952) );
inv1 gate1440( .a(N4832), .O(N5953) );
nand2 gate1441( .a(N4835), .b(N1936), .O(N5954) );
inv1 gate1442( .a(N4835), .O(N5955) );
nand2 gate1443( .a(N4838), .b(N1937), .O(N5956) );
inv1 gate1444( .a(N4838), .O(N5957) );
nand2 gate1445( .a(N4841), .b(N1938), .O(N5958) );
inv1 gate1446( .a(N4841), .O(N5959) );
and2 gate1447( .a(N2674), .b(N4769), .O(N5960) );
inv1 gate1448( .a(N4844), .O(N5966) );
nand2 gate1449( .a(N4847), .b(N1939), .O(N5967) );
inv1 gate1450( .a(N4847), .O(N5968) );
nand2 gate1451( .a(N4850), .b(N1940), .O(N5969) );
inv1 gate1452( .a(N4850), .O(N5970) );
nand2 gate1453( .a(N4853), .b(N1941), .O(N5971) );
inv1 gate1454( .a(N4853), .O(N5972) );
nand2 gate1455( .a(N4856), .b(N1942), .O(N5973) );
inv1 gate1456( .a(N4856), .O(N5974) );
nand2 gate1457( .a(N4859), .b(N1943), .O(N5975) );
inv1 gate1458( .a(N4859), .O(N5976) );
nand2 gate1459( .a(N4862), .b(N1944), .O(N5977) );
inv1 gate1460( .a(N4862), .O(N5978) );
nand2 gate1461( .a(N4865), .b(N1945), .O(N5979) );
inv1 gate1462( .a(N4865), .O(N5980) );
and2 gate1463( .a(N2674), .b(N4769), .O(N5981) );
nand2 gate1464( .a(N4868), .b(N1946), .O(N5989) );
inv1 gate1465( .a(N4868), .O(N5990) );
nand2 gate1466( .a(N5283), .b(N5284), .O(N5991) );
nand2 gate1467( .a(N5285), .b(N5286), .O(N5996) );
nand2 gate1468( .a(N5287), .b(N5288), .O(N6000) );
nand2 gate1469( .a(N5289), .b(N5290), .O(N6003) );
nand2 gate1470( .a(N5291), .b(N5292), .O(N6009) );
nand2 gate1471( .a(N5293), .b(N5294), .O(N6014) );
nand2 gate1472( .a(N5295), .b(N5296), .O(N6018) );
nand2 gate1473( .a(N5297), .b(N5298), .O(N6021) );
nand2 gate1474( .a(N5299), .b(N5300), .O(N6022) );
inv1 gate1475( .a(N4874), .O(N6023) );
nand2 gate1476( .a(N4874), .b(N4629), .O(N6024) );
inv1 gate1477( .a(N4877), .O(N6025) );
nand2 gate1478( .a(N4877), .b(N4631), .O(N6026) );
inv1 gate1479( .a(N4880), .O(N6027) );
nand2 gate1480( .a(N4880), .b(N4633), .O(N6028) );
inv1 gate1481( .a(N4883), .O(N6029) );
nand2 gate1482( .a(N4883), .b(N4636), .O(N6030) );
inv1 gate1483( .a(N4886), .O(N6031) );
inv1 gate1484( .a(N4889), .O(N6032) );
inv1 gate1485( .a(N4892), .O(N6033) );
inv1 gate1486( .a(N4895), .O(N6034) );
inv1 gate1487( .a(N4898), .O(N6035) );
inv1 gate1488( .a(N4901), .O(N6036) );
inv1 gate1489( .a(N4904), .O(N6037) );
nand2 gate1490( .a(N4904), .b(N4642), .O(N6038) );
inv1 gate1491( .a(N4907), .O(N6039) );
inv1 gate1492( .a(N4910), .O(N6040) );
nand2 gate1493( .a(N5314), .b(N5315), .O(N6041) );
inv1 gate( .a(N5316),.O(N5316_NOT) );
inv1 gate( .a(N5317),.O(N5317_NOT));
and2 gate( .a(N5316_NOT), .b(p293), .O(EX731) );
and2 gate( .a(N5317_NOT), .b(EX731), .O(EX732) );
and2 gate( .a(N5316), .b(p294), .O(EX733) );
and2 gate( .a(N5317_NOT), .b(EX733), .O(EX734) );
and2 gate( .a(N5316_NOT), .b(p295), .O(EX735) );
and2 gate( .a(N5317), .b(EX735), .O(EX736) );
and2 gate( .a(N5316), .b(p296), .O(EX737) );
and2 gate( .a(N5317), .b(EX737), .O(EX738) );
or2  gate( .a(EX732), .b(EX734), .O(EX739) );
or2  gate( .a(EX736), .b(EX739), .O(EX740) );
or2  gate( .a(EX738), .b(EX740), .O(N6047) );
nand2 gate1495( .a(N5318), .b(N5319), .O(N6052) );
inv1 gate( .a(N5320),.O(N5320_NOT) );
inv1 gate( .a(N5321),.O(N5321_NOT));
and2 gate( .a(N5320_NOT), .b(p297), .O(EX741) );
and2 gate( .a(N5321_NOT), .b(EX741), .O(EX742) );
and2 gate( .a(N5320), .b(p298), .O(EX743) );
and2 gate( .a(N5321_NOT), .b(EX743), .O(EX744) );
and2 gate( .a(N5320_NOT), .b(p299), .O(EX745) );
and2 gate( .a(N5321), .b(EX745), .O(EX746) );
and2 gate( .a(N5320), .b(p300), .O(EX747) );
and2 gate( .a(N5321), .b(EX747), .O(EX748) );
or2  gate( .a(EX742), .b(EX744), .O(EX749) );
or2  gate( .a(EX746), .b(EX749), .O(EX750) );
or2  gate( .a(EX748), .b(EX750), .O(N6056) );
nand2 gate1497( .a(N5322), .b(N5323), .O(N6059) );
nand2 gate1498( .a(N4913), .b(N1968), .O(N6060) );
inv1 gate1499( .a(N4913), .O(N6061) );
nand2 gate1500( .a(N4916), .b(N1969), .O(N6062) );
inv1 gate1501( .a(N4916), .O(N6063) );
nand2 gate1502( .a(N4919), .b(N1970), .O(N6064) );
inv1 gate1503( .a(N4919), .O(N6065) );
nand2 gate1504( .a(N4922), .b(N1971), .O(N6066) );
inv1 gate1505( .a(N4922), .O(N6067) );
nand2 gate1506( .a(N4925), .b(N1972), .O(N6068) );
inv1 gate1507( .a(N4925), .O(N6069) );
inv1 gate( .a(N4928),.O(N4928_NOT) );
inv1 gate( .a(N1973),.O(N1973_NOT));
and2 gate( .a(N4928_NOT), .b(p301), .O(EX751) );
and2 gate( .a(N1973_NOT), .b(EX751), .O(EX752) );
and2 gate( .a(N4928), .b(p302), .O(EX753) );
and2 gate( .a(N1973_NOT), .b(EX753), .O(EX754) );
and2 gate( .a(N4928_NOT), .b(p303), .O(EX755) );
and2 gate( .a(N1973), .b(EX755), .O(EX756) );
and2 gate( .a(N4928), .b(p304), .O(EX757) );
and2 gate( .a(N1973), .b(EX757), .O(EX758) );
or2  gate( .a(EX752), .b(EX754), .O(EX759) );
or2  gate( .a(EX756), .b(EX759), .O(EX760) );
or2  gate( .a(EX758), .b(EX760), .O(N6070) );
inv1 gate1509( .a(N4928), .O(N6071) );
nand2 gate1510( .a(N4931), .b(N1974), .O(N6072) );
inv1 gate1511( .a(N4931), .O(N6073) );
nand2 gate1512( .a(N4934), .b(N1975), .O(N6074) );
inv1 gate1513( .a(N4934), .O(N6075) );
nand2 gate1514( .a(N4937), .b(N1976), .O(N6076) );
inv1 gate1515( .a(N4937), .O(N6077) );
inv1 gate1516( .a(N4940), .O(N6078) );
nand2 gate1517( .a(N5363), .b(N4694), .O(N6079) );
nand2 gate1518( .a(N5364), .b(N5365), .O(N6083) );
nand2 gate1519( .a(N5366), .b(N5367), .O(N6087) );
inv1 gate1520( .a(N4943), .O(N6090) );
inv1 gate( .a(N4943),.O(N4943_NOT) );
inv1 gate( .a(N4699),.O(N4699_NOT));
and2 gate( .a(N4943_NOT), .b(p305), .O(EX761) );
and2 gate( .a(N4699_NOT), .b(EX761), .O(EX762) );
and2 gate( .a(N4943), .b(p306), .O(EX763) );
and2 gate( .a(N4699_NOT), .b(EX763), .O(EX764) );
and2 gate( .a(N4943_NOT), .b(p307), .O(EX765) );
and2 gate( .a(N4699), .b(EX765), .O(EX766) );
and2 gate( .a(N4943), .b(p308), .O(EX767) );
and2 gate( .a(N4699), .b(EX767), .O(EX768) );
or2  gate( .a(EX762), .b(EX764), .O(EX769) );
or2  gate( .a(EX766), .b(EX769), .O(EX770) );
or2  gate( .a(EX768), .b(EX770), .O(N6091) );
inv1 gate1522( .a(N4946), .O(N6092) );
inv1 gate1523( .a(N4949), .O(N6093) );
inv1 gate1524( .a(N4952), .O(N6094) );
inv1 gate1525( .a(N4955), .O(N6095) );
inv1 gate1526( .a(N4970), .O(N6096) );
nand2 gate1527( .a(N4970), .b(N4700), .O(N6097) );
inv1 gate1528( .a(N4973), .O(N6098) );
inv1 gate1529( .a(N4976), .O(N6099) );
inv1 gate1530( .a(N4979), .O(N6100) );
inv1 gate1531( .a(N4982), .O(N6101) );
inv1 gate1532( .a(N4997), .O(N6102) );
nand2 gate1533( .a(N5000), .b(N2015), .O(N6103) );
inv1 gate1534( .a(N5000), .O(N6104) );
nand2 gate1535( .a(N5003), .b(N2016), .O(N6105) );
inv1 gate1536( .a(N5003), .O(N6106) );
nand2 gate1537( .a(N5006), .b(N2017), .O(N6107) );
inv1 gate1538( .a(N5006), .O(N6108) );
nand2 gate1539( .a(N5009), .b(N2018), .O(N6109) );
inv1 gate1540( .a(N5009), .O(N6110) );
nand2 gate1541( .a(N5012), .b(N2019), .O(N6111) );
inv1 gate1542( .a(N5012), .O(N6112) );
nand2 gate1543( .a(N5015), .b(N2020), .O(N6113) );
inv1 gate1544( .a(N5015), .O(N6114) );
nand2 gate1545( .a(N5018), .b(N2021), .O(N6115) );
inv1 gate1546( .a(N5018), .O(N6116) );
nand2 gate1547( .a(N5021), .b(N2022), .O(N6117) );
inv1 gate1548( .a(N5021), .O(N6118) );
nand2 gate1549( .a(N5024), .b(N2023), .O(N6119) );
inv1 gate1550( .a(N5024), .O(N6120) );
inv1 gate1551( .a(N5033), .O(N6121) );
nand2 gate1552( .a(N5033), .b(N4743), .O(N6122) );
inv1 gate1553( .a(N5036), .O(N6123) );
inv1 gate1554( .a(N5039), .O(N6124) );
nand2 gate1555( .a(N5042), .b(N4744), .O(N6125) );
inv1 gate1556( .a(N5042), .O(N6126) );
nand2 gate1557( .a(N5425), .b(N4746), .O(N6127) );
nand2 gate1558( .a(N5426), .b(N5427), .O(N6131) );
inv1 gate1559( .a(N5049), .O(N6135) );
inv1 gate( .a(N5049),.O(N5049_NOT) );
inv1 gate( .a(N4749),.O(N4749_NOT));
and2 gate( .a(N5049_NOT), .b(p309), .O(EX771) );
and2 gate( .a(N4749_NOT), .b(EX771), .O(EX772) );
and2 gate( .a(N5049), .b(p310), .O(EX773) );
and2 gate( .a(N4749_NOT), .b(EX773), .O(EX774) );
and2 gate( .a(N5049_NOT), .b(p311), .O(EX775) );
and2 gate( .a(N4749), .b(EX775), .O(EX776) );
and2 gate( .a(N5049), .b(p312), .O(EX777) );
and2 gate( .a(N4749), .b(EX777), .O(EX778) );
or2  gate( .a(EX772), .b(EX774), .O(EX779) );
or2  gate( .a(EX776), .b(EX779), .O(EX780) );
or2  gate( .a(EX778), .b(EX780), .O(N6136) );
nand2 gate1561( .a(N5429), .b(N4751), .O(N6137) );
nand2 gate1562( .a(N5430), .b(N5431), .O(N6141) );
nand2 gate1563( .a(N5432), .b(N5433), .O(N6145) );
inv1 gate1564( .a(N5068), .O(N6148) );
inv1 gate1565( .a(N5071), .O(N6149) );
inv1 gate1566( .a(N5074), .O(N6150) );
inv1 gate1567( .a(N5077), .O(N6151) );
inv1 gate1568( .a(N5080), .O(N6152) );
inv1 gate1569( .a(N5083), .O(N6153) );
inv1 gate1570( .a(N5086), .O(N6154) );
inv1 gate1571( .a(N5089), .O(N6155) );
inv1 gate1572( .a(N5092), .O(N6156) );
nand2 gate1573( .a(N5092), .b(N4761), .O(N6157) );
inv1 gate1574( .a(N5095), .O(N6158) );
nand2 gate1575( .a(N5095), .b(N4763), .O(N6159) );
inv1 gate1576( .a(N5098), .O(N6160) );
nand2 gate1577( .a(N5098), .b(N4765), .O(N6161) );
inv1 gate1578( .a(N5101), .O(N6162) );
inv1 gate1579( .a(N5104), .O(N6163) );
nand2 gate1580( .a(N5107), .b(N4768), .O(N6164) );
inv1 gate1581( .a(N5107), .O(N6165) );
nand2 gate1582( .a(N5451), .b(N4776), .O(N6166) );
nand2 gate1583( .a(N5452), .b(N5453), .O(N6170) );
nand2 gate1584( .a(N5454), .b(N5455), .O(N6174) );
nand2 gate1585( .a(N5456), .b(N5457), .O(N6177) );
inv1 gate1586( .a(N5114), .O(N6181) );
inv1 gate1587( .a(N5117), .O(N6182) );
inv1 gate1588( .a(N5120), .O(N6183) );
inv1 gate1589( .a(N5123), .O(N6184) );
inv1 gate1590( .a(N5138), .O(N6185) );
nand2 gate1591( .a(N5138), .b(N4783), .O(N6186) );
inv1 gate1592( .a(N5141), .O(N6187) );
inv1 gate1593( .a(N5144), .O(N6188) );
inv1 gate1594( .a(N5147), .O(N6189) );
inv1 gate1595( .a(N5150), .O(N6190) );
inv1 gate1596( .a(N4784), .O(N6191) );
nand2 gate1597( .a(N4784), .b(N2230), .O(N6192) );
inv1 gate1598( .a(N4790), .O(N6193) );
nand2 gate1599( .a(N4790), .b(N2765), .O(N6194) );
inv1 gate1600( .a(N4796), .O(N6195) );
nand2 gate1601( .a(N5476), .b(N5477), .O(N6196) );
nand2 gate1602( .a(N5474), .b(N5475), .O(N6199) );
inv1 gate1603( .a(N4810), .O(N6202) );
inv1 gate1604( .a(N4814), .O(N6203) );
buf1 gate1605( .a(N4769), .O(N6204) );
buf1 gate1606( .a(N4555), .O(N6207) );
buf1 gate1607( .a(N4769), .O(N6210) );
inv1 gate1608( .a(N4871), .O(N6213) );
buf1 gate1609( .a(N4586), .O(N6214) );
nor2 gate1610( .a(N2674), .b(N4769), .O(N6217) );
buf1 gate1611( .a(N4667), .O(N6220) );
inv1 gate1612( .a(N4958), .O(N6223) );
inv1 gate1613( .a(N4961), .O(N6224) );
inv1 gate1614( .a(N4964), .O(N6225) );
inv1 gate1615( .a(N4967), .O(N6226) );
inv1 gate1616( .a(N4985), .O(N6227) );
inv1 gate1617( .a(N4988), .O(N6228) );
inv1 gate1618( .a(N4991), .O(N6229) );
inv1 gate1619( .a(N4994), .O(N6230) );
inv1 gate1620( .a(N5027), .O(N6231) );
buf1 gate1621( .a(N4711), .O(N6232) );
inv1 gate1622( .a(N5030), .O(N6235) );
buf1 gate1623( .a(N4735), .O(N6236) );
inv1 gate1624( .a(N5052), .O(N6239) );
inv1 gate1625( .a(N5055), .O(N6240) );
inv1 gate1626( .a(N5058), .O(N6241) );
inv1 gate1627( .a(N5061), .O(N6242) );
nand2 gate1628( .a(N5573), .b(N5574), .O(N6243) );
nand2 gate1629( .a(N5571), .b(N5572), .O(N6246) );
nand2 gate1630( .a(N5586), .b(N5587), .O(N6249) );
nand2 gate1631( .a(N5584), .b(N5585), .O(N6252) );
inv1 gate1632( .a(N5126), .O(N6255) );
inv1 gate1633( .a(N5129), .O(N6256) );
inv1 gate1634( .a(N5132), .O(N6257) );
inv1 gate1635( .a(N5135), .O(N6258) );
inv1 gate1636( .a(N5153), .O(N6259) );
inv1 gate1637( .a(N5156), .O(N6260) );
inv1 gate1638( .a(N5159), .O(N6261) );
inv1 gate1639( .a(N5162), .O(N6262) );
nand2 gate1640( .a(N5604), .b(N5605), .O(N6263) );
nand2 gate1641( .a(N5602), .b(N5603), .O(N6266) );
nand2 gate1642( .a(N1380), .b(N5945), .O(N6540) );
nand2 gate1643( .a(N1383), .b(N5947), .O(N6541) );
nand2 gate1644( .a(N1386), .b(N5949), .O(N6542) );
nand2 gate1645( .a(N1389), .b(N5951), .O(N6543) );
nand2 gate1646( .a(N1392), .b(N5953), .O(N6544) );
nand2 gate1647( .a(N1395), .b(N5955), .O(N6545) );
inv1 gate( .a(N1398),.O(N1398_NOT) );
inv1 gate( .a(N5957),.O(N5957_NOT));
and2 gate( .a(N1398_NOT), .b(p313), .O(EX781) );
and2 gate( .a(N5957_NOT), .b(EX781), .O(EX782) );
and2 gate( .a(N1398), .b(p314), .O(EX783) );
and2 gate( .a(N5957_NOT), .b(EX783), .O(EX784) );
and2 gate( .a(N1398_NOT), .b(p315), .O(EX785) );
and2 gate( .a(N5957), .b(EX785), .O(EX786) );
and2 gate( .a(N1398), .b(p316), .O(EX787) );
and2 gate( .a(N5957), .b(EX787), .O(EX788) );
or2  gate( .a(EX782), .b(EX784), .O(EX789) );
or2  gate( .a(EX786), .b(EX789), .O(EX790) );
or2  gate( .a(EX788), .b(EX790), .O(N6546) );
nand2 gate1649( .a(N1401), .b(N5959), .O(N6547) );
nand2 gate1650( .a(N1404), .b(N5968), .O(N6555) );
nand2 gate1651( .a(N1407), .b(N5970), .O(N6556) );
nand2 gate1652( .a(N1410), .b(N5972), .O(N6557) );
nand2 gate1653( .a(N1413), .b(N5974), .O(N6558) );
nand2 gate1654( .a(N1416), .b(N5976), .O(N6559) );
nand2 gate1655( .a(N1419), .b(N5978), .O(N6560) );
nand2 gate1656( .a(N1422), .b(N5980), .O(N6561) );
nand2 gate1657( .a(N1425), .b(N5990), .O(N6569) );
nand2 gate1658( .a(N3721), .b(N6023), .O(N6594) );
nand2 gate1659( .a(N3724), .b(N6025), .O(N6595) );
nand2 gate1660( .a(N3727), .b(N6027), .O(N6596) );
nand2 gate1661( .a(N3730), .b(N6029), .O(N6597) );
inv1 gate( .a(N4889),.O(N4889_NOT) );
inv1 gate( .a(N6031),.O(N6031_NOT));
and2 gate( .a(N4889_NOT), .b(p317), .O(EX791) );
and2 gate( .a(N6031_NOT), .b(EX791), .O(EX792) );
and2 gate( .a(N4889), .b(p318), .O(EX793) );
and2 gate( .a(N6031_NOT), .b(EX793), .O(EX794) );
and2 gate( .a(N4889_NOT), .b(p319), .O(EX795) );
and2 gate( .a(N6031), .b(EX795), .O(EX796) );
and2 gate( .a(N4889), .b(p320), .O(EX797) );
and2 gate( .a(N6031), .b(EX797), .O(EX798) );
or2  gate( .a(EX792), .b(EX794), .O(EX799) );
or2  gate( .a(EX796), .b(EX799), .O(EX800) );
or2  gate( .a(EX798), .b(EX800), .O(N6598) );
nand2 gate1663( .a(N4886), .b(N6032), .O(N6599) );
nand2 gate1664( .a(N4895), .b(N6033), .O(N6600) );
nand2 gate1665( .a(N4892), .b(N6034), .O(N6601) );
nand2 gate1666( .a(N4901), .b(N6035), .O(N6602) );
nand2 gate1667( .a(N4898), .b(N6036), .O(N6603) );
nand2 gate1668( .a(N3733), .b(N6037), .O(N6604) );
nand2 gate1669( .a(N4910), .b(N6039), .O(N6605) );
nand2 gate1670( .a(N4907), .b(N6040), .O(N6606) );
inv1 gate( .a(N1434),.O(N1434_NOT) );
inv1 gate( .a(N6061),.O(N6061_NOT));
and2 gate( .a(N1434_NOT), .b(p321), .O(EX801) );
and2 gate( .a(N6061_NOT), .b(EX801), .O(EX802) );
and2 gate( .a(N1434), .b(p322), .O(EX803) );
and2 gate( .a(N6061_NOT), .b(EX803), .O(EX804) );
and2 gate( .a(N1434_NOT), .b(p323), .O(EX805) );
and2 gate( .a(N6061), .b(EX805), .O(EX806) );
and2 gate( .a(N1434), .b(p324), .O(EX807) );
and2 gate( .a(N6061), .b(EX807), .O(EX808) );
or2  gate( .a(EX802), .b(EX804), .O(EX809) );
or2  gate( .a(EX806), .b(EX809), .O(EX810) );
or2  gate( .a(EX808), .b(EX810), .O(N6621) );
nand2 gate1672( .a(N1437), .b(N6063), .O(N6622) );
nand2 gate1673( .a(N1440), .b(N6065), .O(N6623) );
nand2 gate1674( .a(N1443), .b(N6067), .O(N6624) );
nand2 gate1675( .a(N1446), .b(N6069), .O(N6625) );
nand2 gate1676( .a(N1449), .b(N6071), .O(N6626) );
nand2 gate1677( .a(N1452), .b(N6073), .O(N6627) );
nand2 gate1678( .a(N1455), .b(N6075), .O(N6628) );
nand2 gate1679( .a(N1458), .b(N6077), .O(N6629) );
nand2 gate1680( .a(N3783), .b(N6090), .O(N6639) );
nand2 gate1681( .a(N4949), .b(N6092), .O(N6640) );
nand2 gate1682( .a(N4946), .b(N6093), .O(N6641) );
nand2 gate1683( .a(N4955), .b(N6094), .O(N6642) );
nand2 gate1684( .a(N4952), .b(N6095), .O(N6643) );
nand2 gate1685( .a(N3786), .b(N6096), .O(N6644) );
nand2 gate1686( .a(N4976), .b(N6098), .O(N6645) );
nand2 gate1687( .a(N4973), .b(N6099), .O(N6646) );
nand2 gate1688( .a(N4982), .b(N6100), .O(N6647) );
nand2 gate1689( .a(N4979), .b(N6101), .O(N6648) );
nand2 gate1690( .a(N1461), .b(N6104), .O(N6649) );
nand2 gate1691( .a(N1464), .b(N6106), .O(N6650) );
nand2 gate1692( .a(N1467), .b(N6108), .O(N6651) );
nand2 gate1693( .a(N1470), .b(N6110), .O(N6652) );
nand2 gate1694( .a(N1473), .b(N6112), .O(N6653) );
nand2 gate1695( .a(N1476), .b(N6114), .O(N6654) );
nand2 gate1696( .a(N1479), .b(N6116), .O(N6655) );
nand2 gate1697( .a(N1482), .b(N6118), .O(N6656) );
nand2 gate1698( .a(N1485), .b(N6120), .O(N6657) );
nand2 gate1699( .a(N3789), .b(N6121), .O(N6658) );
nand2 gate1700( .a(N5039), .b(N6123), .O(N6659) );
nand2 gate1701( .a(N5036), .b(N6124), .O(N6660) );
nand2 gate1702( .a(N3792), .b(N6126), .O(N6661) );
nand2 gate1703( .a(N3816), .b(N6135), .O(N6668) );
nand2 gate1704( .a(N5071), .b(N6148), .O(N6677) );
nand2 gate1705( .a(N5068), .b(N6149), .O(N6678) );
nand2 gate1706( .a(N5077), .b(N6150), .O(N6679) );
nand2 gate1707( .a(N5074), .b(N6151), .O(N6680) );
nand2 gate1708( .a(N5083), .b(N6152), .O(N6681) );
nand2 gate1709( .a(N5080), .b(N6153), .O(N6682) );
nand2 gate1710( .a(N5089), .b(N6154), .O(N6683) );
nand2 gate1711( .a(N5086), .b(N6155), .O(N6684) );
nand2 gate1712( .a(N3846), .b(N6156), .O(N6685) );
nand2 gate1713( .a(N3849), .b(N6158), .O(N6686) );
nand2 gate1714( .a(N3852), .b(N6160), .O(N6687) );
nand2 gate1715( .a(N5104), .b(N6162), .O(N6688) );
nand2 gate1716( .a(N5101), .b(N6163), .O(N6689) );
nand2 gate1717( .a(N3855), .b(N6165), .O(N6690) );
inv1 gate( .a(N5117),.O(N5117_NOT) );
inv1 gate( .a(N6181),.O(N6181_NOT));
and2 gate( .a(N5117_NOT), .b(p325), .O(EX811) );
and2 gate( .a(N6181_NOT), .b(EX811), .O(EX812) );
and2 gate( .a(N5117), .b(p326), .O(EX813) );
and2 gate( .a(N6181_NOT), .b(EX813), .O(EX814) );
and2 gate( .a(N5117_NOT), .b(p327), .O(EX815) );
and2 gate( .a(N6181), .b(EX815), .O(EX816) );
and2 gate( .a(N5117), .b(p328), .O(EX817) );
and2 gate( .a(N6181), .b(EX817), .O(EX818) );
or2  gate( .a(EX812), .b(EX814), .O(EX819) );
or2  gate( .a(EX816), .b(EX819), .O(EX820) );
or2  gate( .a(EX818), .b(EX820), .O(N6702) );
nand2 gate1719( .a(N5114), .b(N6182), .O(N6703) );
nand2 gate1720( .a(N5123), .b(N6183), .O(N6704) );
nand2 gate1721( .a(N5120), .b(N6184), .O(N6705) );
nand2 gate1722( .a(N3891), .b(N6185), .O(N6706) );
inv1 gate( .a(N5144),.O(N5144_NOT) );
inv1 gate( .a(N6187),.O(N6187_NOT));
and2 gate( .a(N5144_NOT), .b(p329), .O(EX821) );
and2 gate( .a(N6187_NOT), .b(EX821), .O(EX822) );
and2 gate( .a(N5144), .b(p330), .O(EX823) );
and2 gate( .a(N6187_NOT), .b(EX823), .O(EX824) );
and2 gate( .a(N5144_NOT), .b(p331), .O(EX825) );
and2 gate( .a(N6187), .b(EX825), .O(EX826) );
and2 gate( .a(N5144), .b(p332), .O(EX827) );
and2 gate( .a(N6187), .b(EX827), .O(EX828) );
or2  gate( .a(EX822), .b(EX824), .O(EX829) );
or2  gate( .a(EX826), .b(EX829), .O(EX830) );
or2  gate( .a(EX828), .b(EX830), .O(N6707) );
nand2 gate1724( .a(N5141), .b(N6188), .O(N6708) );
nand2 gate1725( .a(N5150), .b(N6189), .O(N6709) );
nand2 gate1726( .a(N5147), .b(N6190), .O(N6710) );
inv1 gate( .a(N1708),.O(N1708_NOT) );
inv1 gate( .a(N6191),.O(N6191_NOT));
and2 gate( .a(N1708_NOT), .b(p333), .O(EX831) );
and2 gate( .a(N6191_NOT), .b(EX831), .O(EX832) );
and2 gate( .a(N1708), .b(p334), .O(EX833) );
and2 gate( .a(N6191_NOT), .b(EX833), .O(EX834) );
and2 gate( .a(N1708_NOT), .b(p335), .O(EX835) );
and2 gate( .a(N6191), .b(EX835), .O(EX836) );
and2 gate( .a(N1708), .b(p336), .O(EX837) );
and2 gate( .a(N6191), .b(EX837), .O(EX838) );
or2  gate( .a(EX832), .b(EX834), .O(EX839) );
or2  gate( .a(EX836), .b(EX839), .O(EX840) );
or2  gate( .a(EX838), .b(EX840), .O(N6711) );
nand2 gate1728( .a(N2231), .b(N6193), .O(N6712) );
nand2 gate1729( .a(N4961), .b(N6223), .O(N6729) );
nand2 gate1730( .a(N4958), .b(N6224), .O(N6730) );
nand2 gate1731( .a(N4967), .b(N6225), .O(N6731) );
nand2 gate1732( .a(N4964), .b(N6226), .O(N6732) );
nand2 gate1733( .a(N4988), .b(N6227), .O(N6733) );
nand2 gate1734( .a(N4985), .b(N6228), .O(N6734) );
nand2 gate1735( .a(N4994), .b(N6229), .O(N6735) );
nand2 gate1736( .a(N4991), .b(N6230), .O(N6736) );
nand2 gate1737( .a(N5055), .b(N6239), .O(N6741) );
nand2 gate1738( .a(N5052), .b(N6240), .O(N6742) );
nand2 gate1739( .a(N5061), .b(N6241), .O(N6743) );
nand2 gate1740( .a(N5058), .b(N6242), .O(N6744) );
nand2 gate1741( .a(N5129), .b(N6255), .O(N6751) );
nand2 gate1742( .a(N5126), .b(N6256), .O(N6752) );
nand2 gate1743( .a(N5135), .b(N6257), .O(N6753) );
nand2 gate1744( .a(N5132), .b(N6258), .O(N6754) );
nand2 gate1745( .a(N5156), .b(N6259), .O(N6755) );
nand2 gate1746( .a(N5153), .b(N6260), .O(N6756) );
nand2 gate1747( .a(N5162), .b(N6261), .O(N6757) );
nand2 gate1748( .a(N5159), .b(N6262), .O(N6758) );
inv1 gate1749( .a(N5892), .O(N6761) );
and5 gate1750( .a(N5683), .b(N5670), .c(N5654), .d(N5640), .e(N5632), .O(N6762) );
and2 gate1751( .a(N5632), .b(N3097), .O(N6766) );
and3 gate1752( .a(N5640), .b(N5632), .c(N3101), .O(N6767) );
and4 gate1753( .a(N5654), .b(N5632), .c(N3107), .d(N5640), .O(N6768) );
and5 gate1754( .a(N5670), .b(N5654), .c(N5632), .d(N3114), .e(N5640), .O(N6769) );
inv1 gate( .a(N5640),.O(N5640_NOT) );
inv1 gate( .a(N3101),.O(N3101_NOT));
and2 gate( .a(N5640_NOT), .b(p337), .O(EX841) );
and2 gate( .a(N3101_NOT), .b(EX841), .O(EX842) );
and2 gate( .a(N5640), .b(p338), .O(EX843) );
and2 gate( .a(N3101_NOT), .b(EX843), .O(EX844) );
and2 gate( .a(N5640_NOT), .b(p339), .O(EX845) );
and2 gate( .a(N3101), .b(EX845), .O(EX846) );
and2 gate( .a(N5640), .b(p340), .O(EX847) );
and2 gate( .a(N3101), .b(EX847), .O(EX848) );
or2  gate( .a(EX842), .b(EX844), .O(EX849) );
or2  gate( .a(EX846), .b(EX849), .O(EX850) );
or2  gate( .a(EX848), .b(EX850), .O(N6770) );
and3 gate1756( .a(N5654), .b(N3107), .c(N5640), .O(N6771) );
and4 gate1757( .a(N5670), .b(N5654), .c(N3114), .d(N5640), .O(N6772) );
and4 gate1758( .a(N5683), .b(N5654), .c(N5640), .d(N5670), .O(N6773) );
and2 gate1759( .a(N5640), .b(N3101), .O(N6774) );
and3 gate1760( .a(N5654), .b(N3107), .c(N5640), .O(N6775) );
and4 gate1761( .a(N5670), .b(N5654), .c(N3114), .d(N5640), .O(N6776) );
inv1 gate( .a(N5654),.O(N5654_NOT) );
inv1 gate( .a(N3107),.O(N3107_NOT));
and2 gate( .a(N5654_NOT), .b(p341), .O(EX851) );
and2 gate( .a(N3107_NOT), .b(EX851), .O(EX852) );
and2 gate( .a(N5654), .b(p342), .O(EX853) );
and2 gate( .a(N3107_NOT), .b(EX853), .O(EX854) );
and2 gate( .a(N5654_NOT), .b(p343), .O(EX855) );
and2 gate( .a(N3107), .b(EX855), .O(EX856) );
and2 gate( .a(N5654), .b(p344), .O(EX857) );
and2 gate( .a(N3107), .b(EX857), .O(EX858) );
or2  gate( .a(EX852), .b(EX854), .O(EX859) );
or2  gate( .a(EX856), .b(EX859), .O(EX860) );
or2  gate( .a(EX858), .b(EX860), .O(N6777) );
and3 gate1763( .a(N5670), .b(N5654), .c(N3114), .O(N6778) );
and3 gate1764( .a(N5683), .b(N5654), .c(N5670), .O(N6779) );
and2 gate1765( .a(N5654), .b(N3107), .O(N6780) );
and3 gate1766( .a(N5670), .b(N5654), .c(N3114), .O(N6781) );
and2 gate1767( .a(N5670), .b(N3114), .O(N6782) );
and2 gate1768( .a(N5683), .b(N5670), .O(N6783) );
and5 gate1769( .a(N5697), .b(N5728), .c(N5707), .d(N5690), .e(N5718), .O(N6784) );
and2 gate1770( .a(N5690), .b(N3137), .O(N6787) );
and3 gate1771( .a(N5697), .b(N5690), .c(N3140), .O(N6788) );
and4 gate1772( .a(N5707), .b(N5690), .c(N3144), .d(N5697), .O(N6789) );
and5 gate1773( .a(N5718), .b(N5707), .c(N5690), .d(N3149), .e(N5697), .O(N6790) );
and2 gate1774( .a(N5697), .b(N3140), .O(N6791) );
and3 gate1775( .a(N5707), .b(N3144), .c(N5697), .O(N6792) );
and4 gate1776( .a(N5718), .b(N5707), .c(N3149), .d(N5697), .O(N6793) );
and2 gate1777( .a(N3144), .b(N5707), .O(N6794) );
and3 gate1778( .a(N5718), .b(N5707), .c(N3149), .O(N6795) );
and2 gate1779( .a(N5718), .b(N3149), .O(N6796) );
inv1 gate1780( .a(N5736), .O(N6797) );
inv1 gate1781( .a(N5740), .O(N6800) );
inv1 gate1782( .a(N5747), .O(N6803) );
inv1 gate1783( .a(N5751), .O(N6806) );
inv1 gate1784( .a(N5758), .O(N6809) );
inv1 gate1785( .a(N5762), .O(N6812) );
buf1 gate1786( .a(N5744), .O(N6815) );
buf1 gate1787( .a(N5744), .O(N6818) );
buf1 gate1788( .a(N5755), .O(N6821) );
buf1 gate1789( .a(N5755), .O(N6824) );
buf1 gate1790( .a(N5766), .O(N6827) );
buf1 gate1791( .a(N5766), .O(N6830) );
and4 gate1792( .a(N5850), .b(N5789), .c(N5778), .d(N5771), .O(N6833) );
and2 gate1793( .a(N5771), .b(N3169), .O(N6836) );
and3 gate1794( .a(N5778), .b(N5771), .c(N3173), .O(N6837) );
and4 gate1795( .a(N5789), .b(N5771), .c(N3178), .d(N5778), .O(N6838) );
and2 gate1796( .a(N5778), .b(N3173), .O(N6839) );
and3 gate1797( .a(N5789), .b(N3178), .c(N5778), .O(N6840) );
and3 gate1798( .a(N5850), .b(N5789), .c(N5778), .O(N6841) );
and2 gate1799( .a(N5778), .b(N3173), .O(N6842) );
and3 gate1800( .a(N5789), .b(N3178), .c(N5778), .O(N6843) );
and2 gate1801( .a(N5789), .b(N3178), .O(N6844) );
and5 gate1802( .a(N5856), .b(N5837), .c(N5821), .d(N5807), .e(N5799), .O(N6845) );
and2 gate1803( .a(N5799), .b(N3185), .O(N6848) );
and3 gate1804( .a(N5807), .b(N5799), .c(N3189), .O(N6849) );
and4 gate1805( .a(N5821), .b(N5799), .c(N3195), .d(N5807), .O(N6850) );
and5 gate1806( .a(N5837), .b(N5821), .c(N5799), .d(N3202), .e(N5807), .O(N6851) );
and2 gate1807( .a(N5807), .b(N3189), .O(N6852) );
and3 gate1808( .a(N5821), .b(N3195), .c(N5807), .O(N6853) );
and4 gate1809( .a(N5837), .b(N5821), .c(N3202), .d(N5807), .O(N6854) );
and4 gate1810( .a(N5856), .b(N5821), .c(N5807), .d(N5837), .O(N6855) );
and2 gate1811( .a(N5807), .b(N3189), .O(N6856) );
and3 gate1812( .a(N5821), .b(N3195), .c(N5807), .O(N6857) );
and4 gate1813( .a(N5837), .b(N5821), .c(N3202), .d(N5807), .O(N6858) );
and2 gate1814( .a(N5821), .b(N3195), .O(N6859) );
and3 gate1815( .a(N5837), .b(N5821), .c(N3202), .O(N6860) );
and3 gate1816( .a(N5856), .b(N5821), .c(N5837), .O(N6861) );
and2 gate1817( .a(N5821), .b(N3195), .O(N6862) );
and3 gate1818( .a(N5837), .b(N5821), .c(N3202), .O(N6863) );
and2 gate1819( .a(N5837), .b(N3202), .O(N6864) );
inv1 gate( .a(N5850),.O(N5850_NOT) );
inv1 gate( .a(N5789),.O(N5789_NOT));
and2 gate( .a(N5850_NOT), .b(p345), .O(EX861) );
and2 gate( .a(N5789_NOT), .b(EX861), .O(EX862) );
and2 gate( .a(N5850), .b(p346), .O(EX863) );
and2 gate( .a(N5789_NOT), .b(EX863), .O(EX864) );
and2 gate( .a(N5850_NOT), .b(p347), .O(EX865) );
and2 gate( .a(N5789), .b(EX865), .O(EX866) );
and2 gate( .a(N5850), .b(p348), .O(EX867) );
and2 gate( .a(N5789), .b(EX867), .O(EX868) );
or2  gate( .a(EX862), .b(EX864), .O(EX869) );
or2  gate( .a(EX866), .b(EX869), .O(EX870) );
or2  gate( .a(EX868), .b(EX870), .O(N6865) );
inv1 gate( .a(N5856),.O(N5856_NOT) );
inv1 gate( .a(N5837),.O(N5837_NOT));
and2 gate( .a(N5856_NOT), .b(p349), .O(EX871) );
and2 gate( .a(N5837_NOT), .b(EX871), .O(EX872) );
and2 gate( .a(N5856), .b(p350), .O(EX873) );
and2 gate( .a(N5837_NOT), .b(EX873), .O(EX874) );
and2 gate( .a(N5856_NOT), .b(p351), .O(EX875) );
and2 gate( .a(N5837), .b(EX875), .O(EX876) );
and2 gate( .a(N5856), .b(p352), .O(EX877) );
and2 gate( .a(N5837), .b(EX877), .O(EX878) );
or2  gate( .a(EX872), .b(EX874), .O(EX879) );
or2  gate( .a(EX876), .b(EX879), .O(EX880) );
or2  gate( .a(EX878), .b(EX880), .O(N6866) );
and4 gate1822( .a(N5870), .b(N5892), .c(N5881), .d(N5863), .O(N6867) );
and2 gate1823( .a(N5863), .b(N3211), .O(N6870) );
and3 gate1824( .a(N5870), .b(N5863), .c(N3215), .O(N6871) );
and4 gate1825( .a(N5881), .b(N5863), .c(N3221), .d(N5870), .O(N6872) );
inv1 gate( .a(N5870),.O(N5870_NOT) );
inv1 gate( .a(N3215),.O(N3215_NOT));
and2 gate( .a(N5870_NOT), .b(p353), .O(EX881) );
and2 gate( .a(N3215_NOT), .b(EX881), .O(EX882) );
and2 gate( .a(N5870), .b(p354), .O(EX883) );
and2 gate( .a(N3215_NOT), .b(EX883), .O(EX884) );
and2 gate( .a(N5870_NOT), .b(p355), .O(EX885) );
and2 gate( .a(N3215), .b(EX885), .O(EX886) );
and2 gate( .a(N5870), .b(p356), .O(EX887) );
and2 gate( .a(N3215), .b(EX887), .O(EX888) );
or2  gate( .a(EX882), .b(EX884), .O(EX889) );
or2  gate( .a(EX886), .b(EX889), .O(EX890) );
or2  gate( .a(EX888), .b(EX890), .O(N6873) );
and3 gate1827( .a(N5881), .b(N3221), .c(N5870), .O(N6874) );
and3 gate1828( .a(N5892), .b(N5881), .c(N5870), .O(N6875) );
and2 gate1829( .a(N5870), .b(N3215), .O(N6876) );
and3 gate1830( .a(N3221), .b(N5881), .c(N5870), .O(N6877) );
and2 gate1831( .a(N5881), .b(N3221), .O(N6878) );
and2 gate1832( .a(N5892), .b(N5881), .O(N6879) );
and2 gate1833( .a(N5881), .b(N3221), .O(N6880) );
and5 gate1834( .a(N5905), .b(N5936), .c(N5915), .d(N5898), .e(N5926), .O(N6881) );
and2 gate1835( .a(N5898), .b(N3229), .O(N6884) );
and3 gate1836( .a(N5905), .b(N5898), .c(N3232), .O(N6885) );
and4 gate1837( .a(N5915), .b(N5898), .c(N3236), .d(N5905), .O(N6886) );
and5 gate1838( .a(N5926), .b(N5915), .c(N5898), .d(N3241), .e(N5905), .O(N6887) );
and2 gate1839( .a(N5905), .b(N3232), .O(N6888) );
and3 gate1840( .a(N5915), .b(N3236), .c(N5905), .O(N6889) );
and4 gate1841( .a(N5926), .b(N5915), .c(N3241), .d(N5905), .O(N6890) );
inv1 gate( .a(N3236),.O(N3236_NOT) );
inv1 gate( .a(N5915),.O(N5915_NOT));
and2 gate( .a(N3236_NOT), .b(p357), .O(EX891) );
and2 gate( .a(N5915_NOT), .b(EX891), .O(EX892) );
and2 gate( .a(N3236), .b(p358), .O(EX893) );
and2 gate( .a(N5915_NOT), .b(EX893), .O(EX894) );
and2 gate( .a(N3236_NOT), .b(p359), .O(EX895) );
and2 gate( .a(N5915), .b(EX895), .O(EX896) );
and2 gate( .a(N3236), .b(p360), .O(EX897) );
and2 gate( .a(N5915), .b(EX897), .O(EX898) );
or2  gate( .a(EX892), .b(EX894), .O(EX899) );
or2  gate( .a(EX896), .b(EX899), .O(EX900) );
or2  gate( .a(EX898), .b(EX900), .O(N6891) );
and3 gate1843( .a(N5926), .b(N5915), .c(N3241), .O(N6892) );
and2 gate1844( .a(N5926), .b(N3241), .O(N6893) );
nand2 gate1845( .a(N5944), .b(N6540), .O(N6894) );
nand2 gate1846( .a(N5946), .b(N6541), .O(N6901) );
nand2 gate1847( .a(N5948), .b(N6542), .O(N6912) );
nand2 gate1848( .a(N5950), .b(N6543), .O(N6923) );
nand2 gate1849( .a(N5952), .b(N6544), .O(N6929) );
nand2 gate1850( .a(N5954), .b(N6545), .O(N6936) );
nand2 gate1851( .a(N5956), .b(N6546), .O(N6946) );
nand2 gate1852( .a(N5958), .b(N6547), .O(N6957) );
nand2 gate1853( .a(N6204), .b(N4575), .O(N6967) );
inv1 gate1854( .a(N6204), .O(N6968) );
inv1 gate1855( .a(N6207), .O(N6969) );
nand2 gate1856( .a(N5967), .b(N6555), .O(N6970) );
nand2 gate1857( .a(N5969), .b(N6556), .O(N6977) );
nand2 gate1858( .a(N5971), .b(N6557), .O(N6988) );
nand2 gate1859( .a(N5973), .b(N6558), .O(N6998) );
nand2 gate1860( .a(N5975), .b(N6559), .O(N7006) );
nand2 gate1861( .a(N5977), .b(N6560), .O(N7020) );
nand2 gate1862( .a(N5979), .b(N6561), .O(N7036) );
nand2 gate1863( .a(N5989), .b(N6569), .O(N7049) );
nand2 gate1864( .a(N6210), .b(N4610), .O(N7055) );
inv1 gate1865( .a(N6210), .O(N7056) );
and4 gate1866( .a(N6021), .b(N6000), .c(N5996), .d(N5991), .O(N7057) );
and2 gate1867( .a(N5991), .b(N3362), .O(N7060) );
and3 gate1868( .a(N5996), .b(N5991), .c(N3363), .O(N7061) );
and4 gate1869( .a(N6000), .b(N5991), .c(N3364), .d(N5996), .O(N7062) );
and5 gate1870( .a(N6022), .b(N6018), .c(N6014), .d(N6009), .e(N6003), .O(N7063) );
and2 gate1871( .a(N6003), .b(N3366), .O(N7064) );
and3 gate1872( .a(N6009), .b(N6003), .c(N3367), .O(N7065) );
and4 gate1873( .a(N6014), .b(N6003), .c(N3368), .d(N6009), .O(N7066) );
and5 gate1874( .a(N6018), .b(N6014), .c(N6003), .d(N3369), .e(N6009), .O(N7067) );
inv1 gate( .a(N6594),.O(N6594_NOT) );
inv1 gate( .a(N6024),.O(N6024_NOT));
and2 gate( .a(N6594_NOT), .b(p361), .O(EX901) );
and2 gate( .a(N6024_NOT), .b(EX901), .O(EX902) );
and2 gate( .a(N6594), .b(p362), .O(EX903) );
and2 gate( .a(N6024_NOT), .b(EX903), .O(EX904) );
and2 gate( .a(N6594_NOT), .b(p363), .O(EX905) );
and2 gate( .a(N6024), .b(EX905), .O(EX906) );
and2 gate( .a(N6594), .b(p364), .O(EX907) );
and2 gate( .a(N6024), .b(EX907), .O(EX908) );
or2  gate( .a(EX902), .b(EX904), .O(EX909) );
or2  gate( .a(EX906), .b(EX909), .O(EX910) );
or2  gate( .a(EX908), .b(EX910), .O(N7068) );
nand2 gate1876( .a(N6595), .b(N6026), .O(N7073) );
nand2 gate1877( .a(N6596), .b(N6028), .O(N7077) );
inv1 gate( .a(N6597),.O(N6597_NOT) );
inv1 gate( .a(N6030),.O(N6030_NOT));
and2 gate( .a(N6597_NOT), .b(p365), .O(EX911) );
and2 gate( .a(N6030_NOT), .b(EX911), .O(EX912) );
and2 gate( .a(N6597), .b(p366), .O(EX913) );
and2 gate( .a(N6030_NOT), .b(EX913), .O(EX914) );
and2 gate( .a(N6597_NOT), .b(p367), .O(EX915) );
and2 gate( .a(N6030), .b(EX915), .O(EX916) );
and2 gate( .a(N6597), .b(p368), .O(EX917) );
and2 gate( .a(N6030), .b(EX917), .O(EX918) );
or2  gate( .a(EX912), .b(EX914), .O(EX919) );
or2  gate( .a(EX916), .b(EX919), .O(EX920) );
or2  gate( .a(EX918), .b(EX920), .O(N7080) );
nand2 gate1879( .a(N6598), .b(N6599), .O(N7086) );
nand2 gate1880( .a(N6600), .b(N6601), .O(N7091) );
nand2 gate1881( .a(N6602), .b(N6603), .O(N7095) );
nand2 gate1882( .a(N6604), .b(N6038), .O(N7098) );
nand2 gate1883( .a(N6605), .b(N6606), .O(N7099) );
and5 gate1884( .a(N6059), .b(N6056), .c(N6052), .d(N6047), .e(N6041), .O(N7100) );
and2 gate1885( .a(N6041), .b(N3371), .O(N7103) );
and3 gate1886( .a(N6047), .b(N6041), .c(N3372), .O(N7104) );
and4 gate1887( .a(N6052), .b(N6041), .c(N3373), .d(N6047), .O(N7105) );
and5 gate1888( .a(N6056), .b(N6052), .c(N6041), .d(N3374), .e(N6047), .O(N7106) );
nand2 gate1889( .a(N6060), .b(N6621), .O(N7107) );
nand2 gate1890( .a(N6062), .b(N6622), .O(N7114) );
nand2 gate1891( .a(N6064), .b(N6623), .O(N7125) );
nand2 gate1892( .a(N6066), .b(N6624), .O(N7136) );
nand2 gate1893( .a(N6068), .b(N6625), .O(N7142) );
nand2 gate1894( .a(N6070), .b(N6626), .O(N7149) );
nand2 gate1895( .a(N6072), .b(N6627), .O(N7159) );
nand2 gate1896( .a(N6074), .b(N6628), .O(N7170) );
nand2 gate1897( .a(N6076), .b(N6629), .O(N7180) );
inv1 gate1898( .a(N6220), .O(N7187) );
inv1 gate1899( .a(N6079), .O(N7188) );
inv1 gate1900( .a(N6083), .O(N7191) );
nand2 gate1901( .a(N6639), .b(N6091), .O(N7194) );
nand2 gate1902( .a(N6640), .b(N6641), .O(N7198) );
nand2 gate1903( .a(N6642), .b(N6643), .O(N7202) );
nand2 gate1904( .a(N6644), .b(N6097), .O(N7205) );
nand2 gate1905( .a(N6645), .b(N6646), .O(N7209) );
nand2 gate1906( .a(N6647), .b(N6648), .O(N7213) );
buf1 gate1907( .a(N6087), .O(N7216) );
buf1 gate1908( .a(N6087), .O(N7219) );
nand2 gate1909( .a(N6103), .b(N6649), .O(N7222) );
inv1 gate( .a(N6105),.O(N6105_NOT) );
inv1 gate( .a(N6650),.O(N6650_NOT));
and2 gate( .a(N6105_NOT), .b(p369), .O(EX921) );
and2 gate( .a(N6650_NOT), .b(EX921), .O(EX922) );
and2 gate( .a(N6105), .b(p370), .O(EX923) );
and2 gate( .a(N6650_NOT), .b(EX923), .O(EX924) );
and2 gate( .a(N6105_NOT), .b(p371), .O(EX925) );
and2 gate( .a(N6650), .b(EX925), .O(EX926) );
and2 gate( .a(N6105), .b(p372), .O(EX927) );
and2 gate( .a(N6650), .b(EX927), .O(EX928) );
or2  gate( .a(EX922), .b(EX924), .O(EX929) );
or2  gate( .a(EX926), .b(EX929), .O(EX930) );
or2  gate( .a(EX928), .b(EX930), .O(N7229) );
nand2 gate1911( .a(N6107), .b(N6651), .O(N7240) );
nand2 gate1912( .a(N6109), .b(N6652), .O(N7250) );
nand2 gate1913( .a(N6111), .b(N6653), .O(N7258) );
nand2 gate1914( .a(N6113), .b(N6654), .O(N7272) );
inv1 gate( .a(N6115),.O(N6115_NOT) );
inv1 gate( .a(N6655),.O(N6655_NOT));
and2 gate( .a(N6115_NOT), .b(p373), .O(EX931) );
and2 gate( .a(N6655_NOT), .b(EX931), .O(EX932) );
and2 gate( .a(N6115), .b(p374), .O(EX933) );
and2 gate( .a(N6655_NOT), .b(EX933), .O(EX934) );
and2 gate( .a(N6115_NOT), .b(p375), .O(EX935) );
and2 gate( .a(N6655), .b(EX935), .O(EX936) );
and2 gate( .a(N6115), .b(p376), .O(EX937) );
and2 gate( .a(N6655), .b(EX937), .O(EX938) );
or2  gate( .a(EX932), .b(EX934), .O(EX939) );
or2  gate( .a(EX936), .b(EX939), .O(EX940) );
or2  gate( .a(EX938), .b(EX940), .O(N7288) );
nand2 gate1916( .a(N6117), .b(N6656), .O(N7301) );
nand2 gate1917( .a(N6119), .b(N6657), .O(N7307) );
nand2 gate1918( .a(N6658), .b(N6122), .O(N7314) );
nand2 gate1919( .a(N6659), .b(N6660), .O(N7318) );
nand2 gate1920( .a(N6125), .b(N6661), .O(N7322) );
inv1 gate1921( .a(N6127), .O(N7325) );
inv1 gate1922( .a(N6131), .O(N7328) );
nand2 gate1923( .a(N6668), .b(N6136), .O(N7331) );
inv1 gate1924( .a(N6137), .O(N7334) );
inv1 gate1925( .a(N6141), .O(N7337) );
buf1 gate1926( .a(N6145), .O(N7340) );
buf1 gate1927( .a(N6145), .O(N7343) );
inv1 gate( .a(N6677),.O(N6677_NOT) );
inv1 gate( .a(N6678),.O(N6678_NOT));
and2 gate( .a(N6677_NOT), .b(p377), .O(EX941) );
and2 gate( .a(N6678_NOT), .b(EX941), .O(EX942) );
and2 gate( .a(N6677), .b(p378), .O(EX943) );
and2 gate( .a(N6678_NOT), .b(EX943), .O(EX944) );
and2 gate( .a(N6677_NOT), .b(p379), .O(EX945) );
and2 gate( .a(N6678), .b(EX945), .O(EX946) );
and2 gate( .a(N6677), .b(p380), .O(EX947) );
and2 gate( .a(N6678), .b(EX947), .O(EX948) );
or2  gate( .a(EX942), .b(EX944), .O(EX949) );
or2  gate( .a(EX946), .b(EX949), .O(EX950) );
or2  gate( .a(EX948), .b(EX950), .O(N7346) );
nand2 gate1929( .a(N6679), .b(N6680), .O(N7351) );
nand2 gate1930( .a(N6681), .b(N6682), .O(N7355) );
nand2 gate1931( .a(N6683), .b(N6684), .O(N7358) );
nand2 gate1932( .a(N6685), .b(N6157), .O(N7364) );
nand2 gate1933( .a(N6686), .b(N6159), .O(N7369) );
nand2 gate1934( .a(N6687), .b(N6161), .O(N7373) );
nand2 gate1935( .a(N6688), .b(N6689), .O(N7376) );
nand2 gate1936( .a(N6164), .b(N6690), .O(N7377) );
inv1 gate1937( .a(N6166), .O(N7378) );
inv1 gate1938( .a(N6170), .O(N7381) );
inv1 gate1939( .a(N6177), .O(N7384) );
nand2 gate1940( .a(N6702), .b(N6703), .O(N7387) );
nand2 gate1941( .a(N6704), .b(N6705), .O(N7391) );
nand2 gate1942( .a(N6706), .b(N6186), .O(N7394) );
nand2 gate1943( .a(N6707), .b(N6708), .O(N7398) );
nand2 gate1944( .a(N6709), .b(N6710), .O(N7402) );
buf1 gate1945( .a(N6174), .O(N7405) );
buf1 gate1946( .a(N6174), .O(N7408) );
buf1 gate1947( .a(N5936), .O(N7411) );
buf1 gate1948( .a(N5898), .O(N7414) );
buf1 gate1949( .a(N5905), .O(N7417) );
buf1 gate1950( .a(N5915), .O(N7420) );
buf1 gate1951( .a(N5926), .O(N7423) );
buf1 gate1952( .a(N5728), .O(N7426) );
buf1 gate1953( .a(N5690), .O(N7429) );
buf1 gate1954( .a(N5697), .O(N7432) );
buf1 gate1955( .a(N5707), .O(N7435) );
buf1 gate1956( .a(N5718), .O(N7438) );
nand2 gate1957( .a(N6192), .b(N6711), .O(N7441) );
inv1 gate( .a(N6194),.O(N6194_NOT) );
inv1 gate( .a(N6712),.O(N6712_NOT));
and2 gate( .a(N6194_NOT), .b(p381), .O(EX951) );
and2 gate( .a(N6712_NOT), .b(EX951), .O(EX952) );
and2 gate( .a(N6194), .b(p382), .O(EX953) );
and2 gate( .a(N6712_NOT), .b(EX953), .O(EX954) );
and2 gate( .a(N6194_NOT), .b(p383), .O(EX955) );
and2 gate( .a(N6712), .b(EX955), .O(EX956) );
and2 gate( .a(N6194), .b(p384), .O(EX957) );
and2 gate( .a(N6712), .b(EX957), .O(EX958) );
or2  gate( .a(EX952), .b(EX954), .O(EX959) );
or2  gate( .a(EX956), .b(EX959), .O(EX960) );
or2  gate( .a(EX958), .b(EX960), .O(N7444) );
buf1 gate1959( .a(N5683), .O(N7447) );
buf1 gate1960( .a(N5670), .O(N7450) );
buf1 gate1961( .a(N5632), .O(N7453) );
buf1 gate1962( .a(N5654), .O(N7456) );
buf1 gate1963( .a(N5640), .O(N7459) );
buf1 gate1964( .a(N5640), .O(N7462) );
buf1 gate1965( .a(N5683), .O(N7465) );
buf1 gate1966( .a(N5670), .O(N7468) );
buf1 gate1967( .a(N5632), .O(N7471) );
buf1 gate1968( .a(N5654), .O(N7474) );
inv1 gate1969( .a(N6196), .O(N7477) );
inv1 gate1970( .a(N6199), .O(N7478) );
buf1 gate1971( .a(N5850), .O(N7479) );
buf1 gate1972( .a(N5789), .O(N7482) );
buf1 gate1973( .a(N5771), .O(N7485) );
buf1 gate1974( .a(N5778), .O(N7488) );
buf1 gate1975( .a(N5850), .O(N7491) );
buf1 gate1976( .a(N5789), .O(N7494) );
buf1 gate1977( .a(N5771), .O(N7497) );
buf1 gate1978( .a(N5778), .O(N7500) );
buf1 gate1979( .a(N5856), .O(N7503) );
buf1 gate1980( .a(N5837), .O(N7506) );
buf1 gate1981( .a(N5799), .O(N7509) );
buf1 gate1982( .a(N5821), .O(N7512) );
buf1 gate1983( .a(N5807), .O(N7515) );
buf1 gate1984( .a(N5807), .O(N7518) );
buf1 gate1985( .a(N5856), .O(N7521) );
buf1 gate1986( .a(N5837), .O(N7524) );
buf1 gate1987( .a(N5799), .O(N7527) );
buf1 gate1988( .a(N5821), .O(N7530) );
buf1 gate1989( .a(N5863), .O(N7533) );
buf1 gate1990( .a(N5863), .O(N7536) );
buf1 gate1991( .a(N5870), .O(N7539) );
buf1 gate1992( .a(N5870), .O(N7542) );
buf1 gate1993( .a(N5881), .O(N7545) );
buf1 gate1994( .a(N5881), .O(N7548) );
inv1 gate1995( .a(N6214), .O(N7551) );
inv1 gate1996( .a(N6217), .O(N7552) );
buf1 gate1997( .a(N5981), .O(N7553) );
inv1 gate1998( .a(N6249), .O(N7556) );
inv1 gate1999( .a(N6252), .O(N7557) );
inv1 gate2000( .a(N6243), .O(N7558) );
inv1 gate2001( .a(N6246), .O(N7559) );
nand2 gate2002( .a(N6731), .b(N6732), .O(N7560) );
nand2 gate2003( .a(N6729), .b(N6730), .O(N7563) );
nand2 gate2004( .a(N6735), .b(N6736), .O(N7566) );
nand2 gate2005( .a(N6733), .b(N6734), .O(N7569) );
inv1 gate2006( .a(N6232), .O(N7572) );
inv1 gate2007( .a(N6236), .O(N7573) );
inv1 gate( .a(N6743),.O(N6743_NOT) );
inv1 gate( .a(N6744),.O(N6744_NOT));
and2 gate( .a(N6743_NOT), .b(p385), .O(EX961) );
and2 gate( .a(N6744_NOT), .b(EX961), .O(EX962) );
and2 gate( .a(N6743), .b(p386), .O(EX963) );
and2 gate( .a(N6744_NOT), .b(EX963), .O(EX964) );
and2 gate( .a(N6743_NOT), .b(p387), .O(EX965) );
and2 gate( .a(N6744), .b(EX965), .O(EX966) );
and2 gate( .a(N6743), .b(p388), .O(EX967) );
and2 gate( .a(N6744), .b(EX967), .O(EX968) );
or2  gate( .a(EX962), .b(EX964), .O(EX969) );
or2  gate( .a(EX966), .b(EX969), .O(EX970) );
or2  gate( .a(EX968), .b(EX970), .O(N7574) );
nand2 gate2009( .a(N6741), .b(N6742), .O(N7577) );
inv1 gate2010( .a(N6263), .O(N7580) );
inv1 gate2011( .a(N6266), .O(N7581) );
nand2 gate2012( .a(N6753), .b(N6754), .O(N7582) );
nand2 gate2013( .a(N6751), .b(N6752), .O(N7585) );
nand2 gate2014( .a(N6757), .b(N6758), .O(N7588) );
nand2 gate2015( .a(N6755), .b(N6756), .O(N7591) );
or5 gate2016( .a(N3096), .b(N6766), .c(N6767), .d(N6768), .e(N6769), .O(N7609) );
inv1 gate( .a(N3107),.O(N3107_NOT) );
inv1 gate( .a(N6782),.O(N6782_NOT));
and2 gate( .a(N3107_NOT), .b(p389), .O(EX971) );
and2 gate( .a(N6782_NOT), .b(EX971), .O(EX972) );
and2 gate( .a(N3107), .b(p390), .O(EX973) );
and2 gate( .a(N6782_NOT), .b(EX973), .O(EX974) );
and2 gate( .a(N3107_NOT), .b(p391), .O(EX975) );
and2 gate( .a(N6782), .b(EX975), .O(EX976) );
and2 gate( .a(N3107), .b(p392), .O(EX977) );
and2 gate( .a(N6782), .b(EX977), .O(EX978) );
or2  gate( .a(EX972), .b(EX974), .O(EX979) );
or2  gate( .a(EX976), .b(EX979), .O(EX980) );
or2  gate( .a(EX978), .b(EX980), .O(N7613) );
or5 gate2018( .a(N3136), .b(N6787), .c(N6788), .d(N6789), .e(N6790), .O(N7620) );
or4 gate2019( .a(N3168), .b(N6836), .c(N6837), .d(N6838), .O(N7649) );
or2 gate2020( .a(N3173), .b(N6844), .O(N7650) );
or5 gate2021( .a(N3184), .b(N6848), .c(N6849), .d(N6850), .e(N6851), .O(N7655) );
or2 gate2022( .a(N3195), .b(N6864), .O(N7659) );
or4 gate2023( .a(N3210), .b(N6870), .c(N6871), .d(N6872), .O(N7668) );
or5 gate2024( .a(N3228), .b(N6884), .c(N6885), .d(N6886), .e(N6887), .O(N7671) );
nand2 gate2025( .a(N3661), .b(N6968), .O(N7744) );
nand2 gate2026( .a(N3664), .b(N7056), .O(N7822) );
or4 gate2027( .a(N3361), .b(N7060), .c(N7061), .d(N7062), .O(N7825) );
or5 gate2028( .a(N3365), .b(N7064), .c(N7065), .d(N7066), .e(N7067), .O(N7826) );
or5 gate2029( .a(N3370), .b(N7103), .c(N7104), .d(N7105), .e(N7106), .O(N7852) );
or4 gate2030( .a(N3101), .b(N6777), .c(N6778), .d(N6779), .O(N8114) );
or5 gate2031( .a(N3097), .b(N6770), .c(N6771), .d(N6772), .e(N6773), .O(N8117) );
nor3 gate2032( .a(N3101), .b(N6780), .c(N6781), .O(N8131) );
nor4 gate2033( .a(N3097), .b(N6774), .c(N6775), .d(N6776), .O(N8134) );
nand2 gate2034( .a(N6199), .b(N7477), .O(N8144) );
nand2 gate2035( .a(N6196), .b(N7478), .O(N8145) );
or4 gate2036( .a(N3169), .b(N6839), .c(N6840), .d(N6841), .O(N8146) );
nor3 gate2037( .a(N3169), .b(N6842), .c(N6843), .O(N8156) );
or4 gate2038( .a(N3189), .b(N6859), .c(N6860), .d(N6861), .O(N8166) );
or5 gate2039( .a(N3185), .b(N6852), .c(N6853), .d(N6854), .e(N6855), .O(N8169) );
nor3 gate2040( .a(N3189), .b(N6862), .c(N6863), .O(N8183) );
nor4 gate2041( .a(N3185), .b(N6856), .c(N6857), .d(N6858), .O(N8186) );
or4 gate2042( .a(N3211), .b(N6873), .c(N6874), .d(N6875), .O(N8196) );
nor3 gate2043( .a(N3211), .b(N6876), .c(N6877), .O(N8200) );
or3 gate2044( .a(N3215), .b(N6878), .c(N6879), .O(N8204) );
nor2 gate2045( .a(N3215), .b(N6880), .O(N8208) );
nand2 gate2046( .a(N6252), .b(N7556), .O(N8216) );
nand2 gate2047( .a(N6249), .b(N7557), .O(N8217) );
nand2 gate2048( .a(N6246), .b(N7558), .O(N8218) );
nand2 gate2049( .a(N6243), .b(N7559), .O(N8219) );
nand2 gate2050( .a(N6266), .b(N7580), .O(N8232) );
nand2 gate2051( .a(N6263), .b(N7581), .O(N8233) );
inv1 gate2052( .a(N7411), .O(N8242) );
inv1 gate2053( .a(N7414), .O(N8243) );
inv1 gate2054( .a(N7417), .O(N8244) );
inv1 gate2055( .a(N7420), .O(N8245) );
inv1 gate2056( .a(N7423), .O(N8246) );
inv1 gate2057( .a(N7426), .O(N8247) );
inv1 gate2058( .a(N7429), .O(N8248) );
inv1 gate2059( .a(N7432), .O(N8249) );
inv1 gate2060( .a(N7435), .O(N8250) );
inv1 gate2061( .a(N7438), .O(N8251) );
inv1 gate2062( .a(N7136), .O(N8252) );
inv1 gate2063( .a(N6923), .O(N8253) );
inv1 gate2064( .a(N6762), .O(N8254) );
inv1 gate2065( .a(N7459), .O(N8260) );
inv1 gate2066( .a(N7462), .O(N8261) );
and2 gate2067( .a(N3122), .b(N6762), .O(N8262) );
and2 gate2068( .a(N3155), .b(N6784), .O(N8269) );
inv1 gate2069( .a(N6815), .O(N8274) );
inv1 gate2070( .a(N6818), .O(N8275) );
inv1 gate2071( .a(N6821), .O(N8276) );
inv1 gate2072( .a(N6824), .O(N8277) );
inv1 gate2073( .a(N6827), .O(N8278) );
inv1 gate2074( .a(N6830), .O(N8279) );
and3 gate2075( .a(N5740), .b(N5736), .c(N6815), .O(N8280) );
and3 gate2076( .a(N6800), .b(N6797), .c(N6818), .O(N8281) );
and3 gate2077( .a(N5751), .b(N5747), .c(N6821), .O(N8282) );
and3 gate2078( .a(N6806), .b(N6803), .c(N6824), .O(N8283) );
and3 gate2079( .a(N5762), .b(N5758), .c(N6827), .O(N8284) );
and3 gate2080( .a(N6812), .b(N6809), .c(N6830), .O(N8285) );
inv1 gate2081( .a(N6845), .O(N8288) );
inv1 gate2082( .a(N7488), .O(N8294) );
inv1 gate2083( .a(N7500), .O(N8295) );
inv1 gate2084( .a(N7515), .O(N8296) );
inv1 gate2085( .a(N7518), .O(N8297) );
inv1 gate( .a(N6833),.O(N6833_NOT) );
inv1 gate( .a(N6845),.O(N6845_NOT));
and2 gate( .a(N6833_NOT), .b(p393), .O(EX981) );
and2 gate( .a(N6845_NOT), .b(EX981), .O(EX982) );
and2 gate( .a(N6833), .b(p394), .O(EX983) );
and2 gate( .a(N6845_NOT), .b(EX983), .O(EX984) );
and2 gate( .a(N6833_NOT), .b(p395), .O(EX985) );
and2 gate( .a(N6845), .b(EX985), .O(EX986) );
and2 gate( .a(N6833), .b(p396), .O(EX987) );
and2 gate( .a(N6845), .b(EX987), .O(EX988) );
or2  gate( .a(EX982), .b(EX984), .O(EX989) );
or2  gate( .a(EX986), .b(EX989), .O(EX990) );
or2  gate( .a(EX988), .b(EX990), .O(N8298) );
and2 gate2087( .a(N6867), .b(N6881), .O(N8307) );
inv1 gate2088( .a(N7533), .O(N8315) );
inv1 gate2089( .a(N7536), .O(N8317) );
inv1 gate2090( .a(N7539), .O(N8319) );
inv1 gate2091( .a(N7542), .O(N8321) );
nand2 gate2092( .a(N7545), .b(N4543), .O(N8322) );
inv1 gate2093( .a(N7545), .O(N8323) );
nand2 gate2094( .a(N7548), .b(N5943), .O(N8324) );
inv1 gate2095( .a(N7548), .O(N8325) );
nand2 gate2096( .a(N6967), .b(N7744), .O(N8326) );
and4 gate2097( .a(N6901), .b(N6923), .c(N6912), .d(N6894), .O(N8333) );
and2 gate2098( .a(N6894), .b(N4545), .O(N8337) );
and3 gate2099( .a(N6901), .b(N6894), .c(N4549), .O(N8338) );
and4 gate2100( .a(N6912), .b(N6894), .c(N4555), .d(N6901), .O(N8339) );
and2 gate2101( .a(N6901), .b(N4549), .O(N8340) );
and3 gate2102( .a(N6912), .b(N4555), .c(N6901), .O(N8341) );
and3 gate2103( .a(N6923), .b(N6912), .c(N6901), .O(N8342) );
and2 gate2104( .a(N6901), .b(N4549), .O(N8343) );
and3 gate2105( .a(N4555), .b(N6912), .c(N6901), .O(N8344) );
and2 gate2106( .a(N6912), .b(N4555), .O(N8345) );
and2 gate2107( .a(N6923), .b(N6912), .O(N8346) );
and2 gate2108( .a(N6912), .b(N4555), .O(N8347) );
and2 gate2109( .a(N6929), .b(N4563), .O(N8348) );
and3 gate2110( .a(N6936), .b(N6929), .c(N4566), .O(N8349) );
and4 gate2111( .a(N6946), .b(N6929), .c(N4570), .d(N6936), .O(N8350) );
and5 gate2112( .a(N6957), .b(N6946), .c(N6929), .d(N5960), .e(N6936), .O(N8351) );
and2 gate2113( .a(N6936), .b(N4566), .O(N8352) );
and3 gate2114( .a(N6946), .b(N4570), .c(N6936), .O(N8353) );
and4 gate2115( .a(N6957), .b(N6946), .c(N5960), .d(N6936), .O(N8354) );
and2 gate2116( .a(N4570), .b(N6946), .O(N8355) );
and3 gate2117( .a(N6957), .b(N6946), .c(N5960), .O(N8356) );
and2 gate2118( .a(N6957), .b(N5960), .O(N8357) );
nand2 gate2119( .a(N7055), .b(N7822), .O(N8358) );
and4 gate2120( .a(N7049), .b(N6988), .c(N6977), .d(N6970), .O(N8365) );
and2 gate2121( .a(N6970), .b(N4577), .O(N8369) );
and3 gate2122( .a(N6977), .b(N6970), .c(N4581), .O(N8370) );
and4 gate2123( .a(N6988), .b(N6970), .c(N4586), .d(N6977), .O(N8371) );
inv1 gate( .a(N6977),.O(N6977_NOT) );
inv1 gate( .a(N4581),.O(N4581_NOT));
and2 gate( .a(N6977_NOT), .b(p397), .O(EX991) );
and2 gate( .a(N4581_NOT), .b(EX991), .O(EX992) );
and2 gate( .a(N6977), .b(p398), .O(EX993) );
and2 gate( .a(N4581_NOT), .b(EX993), .O(EX994) );
and2 gate( .a(N6977_NOT), .b(p399), .O(EX995) );
and2 gate( .a(N4581), .b(EX995), .O(EX996) );
and2 gate( .a(N6977), .b(p400), .O(EX997) );
and2 gate( .a(N4581), .b(EX997), .O(EX998) );
or2  gate( .a(EX992), .b(EX994), .O(EX999) );
or2  gate( .a(EX996), .b(EX999), .O(EX1000) );
or2  gate( .a(EX998), .b(EX1000), .O(N8372) );
and3 gate2125( .a(N6988), .b(N4586), .c(N6977), .O(N8373) );
and3 gate2126( .a(N7049), .b(N6988), .c(N6977), .O(N8374) );
and2 gate2127( .a(N6977), .b(N4581), .O(N8375) );
and3 gate2128( .a(N6988), .b(N4586), .c(N6977), .O(N8376) );
and2 gate2129( .a(N6988), .b(N4586), .O(N8377) );
and2 gate2130( .a(N6998), .b(N4593), .O(N8378) );
and3 gate2131( .a(N7006), .b(N6998), .c(N4597), .O(N8379) );
and4 gate2132( .a(N7020), .b(N6998), .c(N4603), .d(N7006), .O(N8380) );
and5 gate2133( .a(N7036), .b(N7020), .c(N6998), .d(N5981), .e(N7006), .O(N8381) );
and2 gate2134( .a(N7006), .b(N4597), .O(N8382) );
and3 gate2135( .a(N7020), .b(N4603), .c(N7006), .O(N8383) );
and4 gate2136( .a(N7036), .b(N7020), .c(N5981), .d(N7006), .O(N8384) );
and2 gate2137( .a(N7006), .b(N4597), .O(N8385) );
and3 gate2138( .a(N7020), .b(N4603), .c(N7006), .O(N8386) );
and4 gate2139( .a(N7036), .b(N7020), .c(N5981), .d(N7006), .O(N8387) );
and2 gate2140( .a(N7020), .b(N4603), .O(N8388) );
and3 gate2141( .a(N7036), .b(N7020), .c(N5981), .O(N8389) );
and2 gate2142( .a(N7020), .b(N4603), .O(N8390) );
and3 gate2143( .a(N7036), .b(N7020), .c(N5981), .O(N8391) );
and2 gate2144( .a(N7036), .b(N5981), .O(N8392) );
and2 gate2145( .a(N7049), .b(N6988), .O(N8393) );
inv1 gate( .a(N7057),.O(N7057_NOT) );
inv1 gate( .a(N7063),.O(N7063_NOT));
and2 gate( .a(N7057_NOT), .b(p401), .O(EX1001) );
and2 gate( .a(N7063_NOT), .b(EX1001), .O(EX1002) );
and2 gate( .a(N7057), .b(p402), .O(EX1003) );
and2 gate( .a(N7063_NOT), .b(EX1003), .O(EX1004) );
and2 gate( .a(N7057_NOT), .b(p403), .O(EX1005) );
and2 gate( .a(N7063), .b(EX1005), .O(EX1006) );
and2 gate( .a(N7057), .b(p404), .O(EX1007) );
and2 gate( .a(N7063), .b(EX1007), .O(EX1008) );
or2  gate( .a(EX1002), .b(EX1004), .O(EX1009) );
or2  gate( .a(EX1006), .b(EX1009), .O(EX1010) );
or2  gate( .a(EX1008), .b(EX1010), .O(N8394) );
and2 gate2147( .a(N7057), .b(N7826), .O(N8404) );
and4 gate2148( .a(N7098), .b(N7077), .c(N7073), .d(N7068), .O(N8405) );
and2 gate2149( .a(N7068), .b(N4632), .O(N8409) );
and3 gate2150( .a(N7073), .b(N7068), .c(N4634), .O(N8410) );
and4 gate2151( .a(N7077), .b(N7068), .c(N4635), .d(N7073), .O(N8411) );
and5 gate2152( .a(N7099), .b(N7095), .c(N7091), .d(N7086), .e(N7080), .O(N8412) );
and2 gate2153( .a(N7080), .b(N4638), .O(N8415) );
and3 gate2154( .a(N7086), .b(N7080), .c(N4639), .O(N8416) );
and4 gate2155( .a(N7091), .b(N7080), .c(N4640), .d(N7086), .O(N8417) );
and5 gate2156( .a(N7095), .b(N7091), .c(N7080), .d(N4641), .e(N7086), .O(N8418) );
inv1 gate( .a(N3375),.O(N3375_NOT) );
inv1 gate( .a(N7100),.O(N7100_NOT));
and2 gate( .a(N3375_NOT), .b(p405), .O(EX1011) );
and2 gate( .a(N7100_NOT), .b(EX1011), .O(EX1012) );
and2 gate( .a(N3375), .b(p406), .O(EX1013) );
and2 gate( .a(N7100_NOT), .b(EX1013), .O(EX1014) );
and2 gate( .a(N3375_NOT), .b(p407), .O(EX1015) );
and2 gate( .a(N7100), .b(EX1015), .O(EX1016) );
and2 gate( .a(N3375), .b(p408), .O(EX1017) );
and2 gate( .a(N7100), .b(EX1017), .O(EX1018) );
or2  gate( .a(EX1012), .b(EX1014), .O(EX1019) );
or2  gate( .a(EX1016), .b(EX1019), .O(EX1020) );
or2  gate( .a(EX1018), .b(EX1020), .O(N8421) );
and4 gate2158( .a(N7114), .b(N7136), .c(N7125), .d(N7107), .O(N8430) );
and2 gate2159( .a(N7107), .b(N4657), .O(N8433) );
and3 gate2160( .a(N7114), .b(N7107), .c(N4661), .O(N8434) );
and4 gate2161( .a(N7125), .b(N7107), .c(N4667), .d(N7114), .O(N8435) );
and2 gate2162( .a(N7114), .b(N4661), .O(N8436) );
and3 gate2163( .a(N7125), .b(N4667), .c(N7114), .O(N8437) );
and3 gate2164( .a(N7136), .b(N7125), .c(N7114), .O(N8438) );
and2 gate2165( .a(N7114), .b(N4661), .O(N8439) );
and3 gate2166( .a(N4667), .b(N7125), .c(N7114), .O(N8440) );
inv1 gate( .a(N7125),.O(N7125_NOT) );
inv1 gate( .a(N4667),.O(N4667_NOT));
and2 gate( .a(N7125_NOT), .b(p409), .O(EX1021) );
and2 gate( .a(N4667_NOT), .b(EX1021), .O(EX1022) );
and2 gate( .a(N7125), .b(p410), .O(EX1023) );
and2 gate( .a(N4667_NOT), .b(EX1023), .O(EX1024) );
and2 gate( .a(N7125_NOT), .b(p411), .O(EX1025) );
and2 gate( .a(N4667), .b(EX1025), .O(EX1026) );
and2 gate( .a(N7125), .b(p412), .O(EX1027) );
and2 gate( .a(N4667), .b(EX1027), .O(EX1028) );
or2  gate( .a(EX1022), .b(EX1024), .O(EX1029) );
or2  gate( .a(EX1026), .b(EX1029), .O(EX1030) );
or2  gate( .a(EX1028), .b(EX1030), .O(N8441) );
and2 gate2168( .a(N7136), .b(N7125), .O(N8442) );
and2 gate2169( .a(N7125), .b(N4667), .O(N8443) );
and5 gate2170( .a(N7149), .b(N7180), .c(N7159), .d(N7142), .e(N7170), .O(N8444) );
and2 gate2171( .a(N7142), .b(N4675), .O(N8447) );
and3 gate2172( .a(N7149), .b(N7142), .c(N4678), .O(N8448) );
and4 gate2173( .a(N7159), .b(N7142), .c(N4682), .d(N7149), .O(N8449) );
and5 gate2174( .a(N7170), .b(N7159), .c(N7142), .d(N4687), .e(N7149), .O(N8450) );
and2 gate2175( .a(N7149), .b(N4678), .O(N8451) );
and3 gate2176( .a(N7159), .b(N4682), .c(N7149), .O(N8452) );
and4 gate2177( .a(N7170), .b(N7159), .c(N4687), .d(N7149), .O(N8453) );
and2 gate2178( .a(N4682), .b(N7159), .O(N8454) );
and3 gate2179( .a(N7170), .b(N7159), .c(N4687), .O(N8455) );
and2 gate2180( .a(N7170), .b(N4687), .O(N8456) );
inv1 gate2181( .a(N7194), .O(N8457) );
inv1 gate2182( .a(N7198), .O(N8460) );
inv1 gate2183( .a(N7205), .O(N8463) );
inv1 gate2184( .a(N7209), .O(N8466) );
inv1 gate2185( .a(N7216), .O(N8469) );
inv1 gate2186( .a(N7219), .O(N8470) );
buf1 gate2187( .a(N7202), .O(N8471) );
buf1 gate2188( .a(N7202), .O(N8474) );
buf1 gate2189( .a(N7213), .O(N8477) );
buf1 gate2190( .a(N7213), .O(N8480) );
and3 gate2191( .a(N6083), .b(N6079), .c(N7216), .O(N8483) );
and3 gate2192( .a(N7191), .b(N7188), .c(N7219), .O(N8484) );
and4 gate2193( .a(N7301), .b(N7240), .c(N7229), .d(N7222), .O(N8485) );
and2 gate2194( .a(N7222), .b(N4702), .O(N8488) );
and3 gate2195( .a(N7229), .b(N7222), .c(N4706), .O(N8489) );
and4 gate2196( .a(N7240), .b(N7222), .c(N4711), .d(N7229), .O(N8490) );
and2 gate2197( .a(N7229), .b(N4706), .O(N8491) );
and3 gate2198( .a(N7240), .b(N4711), .c(N7229), .O(N8492) );
and3 gate2199( .a(N7301), .b(N7240), .c(N7229), .O(N8493) );
and2 gate2200( .a(N7229), .b(N4706), .O(N8494) );
and3 gate2201( .a(N7240), .b(N4711), .c(N7229), .O(N8495) );
and2 gate2202( .a(N7240), .b(N4711), .O(N8496) );
and5 gate2203( .a(N7307), .b(N7288), .c(N7272), .d(N7258), .e(N7250), .O(N8497) );
and2 gate2204( .a(N7250), .b(N4718), .O(N8500) );
and3 gate2205( .a(N7258), .b(N7250), .c(N4722), .O(N8501) );
and4 gate2206( .a(N7272), .b(N7250), .c(N4728), .d(N7258), .O(N8502) );
and5 gate2207( .a(N7288), .b(N7272), .c(N7250), .d(N4735), .e(N7258), .O(N8503) );
inv1 gate( .a(N7258),.O(N7258_NOT) );
inv1 gate( .a(N4722),.O(N4722_NOT));
and2 gate( .a(N7258_NOT), .b(p413), .O(EX1031) );
and2 gate( .a(N4722_NOT), .b(EX1031), .O(EX1032) );
and2 gate( .a(N7258), .b(p414), .O(EX1033) );
and2 gate( .a(N4722_NOT), .b(EX1033), .O(EX1034) );
and2 gate( .a(N7258_NOT), .b(p415), .O(EX1035) );
and2 gate( .a(N4722), .b(EX1035), .O(EX1036) );
and2 gate( .a(N7258), .b(p416), .O(EX1037) );
and2 gate( .a(N4722), .b(EX1037), .O(EX1038) );
or2  gate( .a(EX1032), .b(EX1034), .O(EX1039) );
or2  gate( .a(EX1036), .b(EX1039), .O(EX1040) );
or2  gate( .a(EX1038), .b(EX1040), .O(N8504) );
and3 gate2209( .a(N7272), .b(N4728), .c(N7258), .O(N8505) );
and4 gate2210( .a(N7288), .b(N7272), .c(N4735), .d(N7258), .O(N8506) );
and4 gate2211( .a(N7307), .b(N7272), .c(N7258), .d(N7288), .O(N8507) );
and2 gate2212( .a(N7258), .b(N4722), .O(N8508) );
and3 gate2213( .a(N7272), .b(N4728), .c(N7258), .O(N8509) );
and4 gate2214( .a(N7288), .b(N7272), .c(N4735), .d(N7258), .O(N8510) );
and2 gate2215( .a(N7272), .b(N4728), .O(N8511) );
and3 gate2216( .a(N7288), .b(N7272), .c(N4735), .O(N8512) );
and3 gate2217( .a(N7307), .b(N7272), .c(N7288), .O(N8513) );
and2 gate2218( .a(N7272), .b(N4728), .O(N8514) );
and3 gate2219( .a(N7288), .b(N7272), .c(N4735), .O(N8515) );
and2 gate2220( .a(N7288), .b(N4735), .O(N8516) );
and2 gate2221( .a(N7301), .b(N7240), .O(N8517) );
inv1 gate( .a(N7307),.O(N7307_NOT) );
inv1 gate( .a(N7288),.O(N7288_NOT));
and2 gate( .a(N7307_NOT), .b(p417), .O(EX1041) );
and2 gate( .a(N7288_NOT), .b(EX1041), .O(EX1042) );
and2 gate( .a(N7307), .b(p418), .O(EX1043) );
and2 gate( .a(N7288_NOT), .b(EX1043), .O(EX1044) );
and2 gate( .a(N7307_NOT), .b(p419), .O(EX1045) );
and2 gate( .a(N7288), .b(EX1045), .O(EX1046) );
and2 gate( .a(N7307), .b(p420), .O(EX1047) );
and2 gate( .a(N7288), .b(EX1047), .O(EX1048) );
or2  gate( .a(EX1042), .b(EX1044), .O(EX1049) );
or2  gate( .a(EX1046), .b(EX1049), .O(EX1050) );
or2  gate( .a(EX1048), .b(EX1050), .O(N8518) );
inv1 gate2223( .a(N7314), .O(N8519) );
inv1 gate2224( .a(N7318), .O(N8522) );
buf1 gate2225( .a(N7322), .O(N8525) );
buf1 gate2226( .a(N7322), .O(N8528) );
buf1 gate2227( .a(N7331), .O(N8531) );
buf1 gate2228( .a(N7331), .O(N8534) );
inv1 gate2229( .a(N7340), .O(N8537) );
inv1 gate2230( .a(N7343), .O(N8538) );
and3 gate2231( .a(N6141), .b(N6137), .c(N7340), .O(N8539) );
and3 gate2232( .a(N7337), .b(N7334), .c(N7343), .O(N8540) );
and4 gate2233( .a(N7376), .b(N7355), .c(N7351), .d(N7346), .O(N8541) );
and2 gate2234( .a(N7346), .b(N4757), .O(N8545) );
and3 gate2235( .a(N7351), .b(N7346), .c(N4758), .O(N8546) );
and4 gate2236( .a(N7355), .b(N7346), .c(N4759), .d(N7351), .O(N8547) );
and5 gate2237( .a(N7377), .b(N7373), .c(N7369), .d(N7364), .e(N7358), .O(N8548) );
and2 gate2238( .a(N7358), .b(N4762), .O(N8551) );
and3 gate2239( .a(N7364), .b(N7358), .c(N4764), .O(N8552) );
and4 gate2240( .a(N7369), .b(N7358), .c(N4766), .d(N7364), .O(N8553) );
and5 gate2241( .a(N7373), .b(N7369), .c(N7358), .d(N4767), .e(N7364), .O(N8554) );
inv1 gate2242( .a(N7387), .O(N8555) );
inv1 gate2243( .a(N7394), .O(N8558) );
inv1 gate2244( .a(N7398), .O(N8561) );
inv1 gate2245( .a(N7405), .O(N8564) );
inv1 gate2246( .a(N7408), .O(N8565) );
buf1 gate2247( .a(N7391), .O(N8566) );
buf1 gate2248( .a(N7391), .O(N8569) );
buf1 gate2249( .a(N7402), .O(N8572) );
buf1 gate2250( .a(N7402), .O(N8575) );
and3 gate2251( .a(N6170), .b(N6166), .c(N7405), .O(N8578) );
and3 gate2252( .a(N7381), .b(N7378), .c(N7408), .O(N8579) );
buf1 gate2253( .a(N7180), .O(N8580) );
buf1 gate2254( .a(N7142), .O(N8583) );
buf1 gate2255( .a(N7149), .O(N8586) );
buf1 gate2256( .a(N7159), .O(N8589) );
buf1 gate2257( .a(N7170), .O(N8592) );
buf1 gate2258( .a(N6929), .O(N8595) );
buf1 gate2259( .a(N6936), .O(N8598) );
buf1 gate2260( .a(N6946), .O(N8601) );
buf1 gate2261( .a(N6957), .O(N8604) );
inv1 gate2262( .a(N7441), .O(N8607) );
nand2 gate2263( .a(N7441), .b(N5469), .O(N8608) );
inv1 gate2264( .a(N7444), .O(N8609) );
nand2 gate2265( .a(N7444), .b(N4793), .O(N8610) );
inv1 gate2266( .a(N7447), .O(N8615) );
inv1 gate2267( .a(N7450), .O(N8616) );
inv1 gate2268( .a(N7453), .O(N8617) );
inv1 gate2269( .a(N7456), .O(N8618) );
inv1 gate2270( .a(N7474), .O(N8619) );
inv1 gate2271( .a(N7465), .O(N8624) );
inv1 gate2272( .a(N7468), .O(N8625) );
inv1 gate2273( .a(N7471), .O(N8626) );
nand2 gate2274( .a(N8144), .b(N8145), .O(N8627) );
inv1 gate2275( .a(N7479), .O(N8632) );
inv1 gate2276( .a(N7482), .O(N8633) );
inv1 gate2277( .a(N7485), .O(N8634) );
inv1 gate2278( .a(N7491), .O(N8637) );
inv1 gate2279( .a(N7494), .O(N8638) );
inv1 gate2280( .a(N7497), .O(N8639) );
inv1 gate2281( .a(N7503), .O(N8644) );
inv1 gate2282( .a(N7506), .O(N8645) );
inv1 gate2283( .a(N7509), .O(N8646) );
inv1 gate2284( .a(N7512), .O(N8647) );
inv1 gate2285( .a(N7530), .O(N8648) );
inv1 gate2286( .a(N7521), .O(N8653) );
inv1 gate2287( .a(N7524), .O(N8654) );
inv1 gate2288( .a(N7527), .O(N8655) );
buf1 gate2289( .a(N6894), .O(N8660) );
buf1 gate2290( .a(N6894), .O(N8663) );
buf1 gate2291( .a(N6901), .O(N8666) );
buf1 gate2292( .a(N6901), .O(N8669) );
buf1 gate2293( .a(N6912), .O(N8672) );
buf1 gate2294( .a(N6912), .O(N8675) );
buf1 gate2295( .a(N7049), .O(N8678) );
buf1 gate2296( .a(N6988), .O(N8681) );
buf1 gate2297( .a(N6970), .O(N8684) );
buf1 gate2298( .a(N6977), .O(N8687) );
buf1 gate2299( .a(N7049), .O(N8690) );
buf1 gate2300( .a(N6988), .O(N8693) );
buf1 gate2301( .a(N6970), .O(N8696) );
buf1 gate2302( .a(N6977), .O(N8699) );
buf1 gate2303( .a(N7036), .O(N8702) );
buf1 gate2304( .a(N6998), .O(N8705) );
buf1 gate2305( .a(N7020), .O(N8708) );
buf1 gate2306( .a(N7006), .O(N8711) );
buf1 gate2307( .a(N7006), .O(N8714) );
inv1 gate2308( .a(N7553), .O(N8717) );
buf1 gate2309( .a(N7036), .O(N8718) );
buf1 gate2310( .a(N6998), .O(N8721) );
buf1 gate2311( .a(N7020), .O(N8724) );
nand2 gate2312( .a(N8216), .b(N8217), .O(N8727) );
nand2 gate2313( .a(N8218), .b(N8219), .O(N8730) );
inv1 gate2314( .a(N7574), .O(N8733) );
inv1 gate2315( .a(N7577), .O(N8734) );
buf1 gate2316( .a(N7107), .O(N8735) );
buf1 gate2317( .a(N7107), .O(N8738) );
buf1 gate2318( .a(N7114), .O(N8741) );
buf1 gate2319( .a(N7114), .O(N8744) );
buf1 gate2320( .a(N7125), .O(N8747) );
buf1 gate2321( .a(N7125), .O(N8750) );
inv1 gate2322( .a(N7560), .O(N8753) );
inv1 gate2323( .a(N7563), .O(N8754) );
inv1 gate2324( .a(N7566), .O(N8755) );
inv1 gate2325( .a(N7569), .O(N8756) );
buf1 gate2326( .a(N7301), .O(N8757) );
buf1 gate2327( .a(N7240), .O(N8760) );
buf1 gate2328( .a(N7222), .O(N8763) );
buf1 gate2329( .a(N7229), .O(N8766) );
buf1 gate2330( .a(N7301), .O(N8769) );
buf1 gate2331( .a(N7240), .O(N8772) );
buf1 gate2332( .a(N7222), .O(N8775) );
buf1 gate2333( .a(N7229), .O(N8778) );
buf1 gate2334( .a(N7307), .O(N8781) );
buf1 gate2335( .a(N7288), .O(N8784) );
buf1 gate2336( .a(N7250), .O(N8787) );
buf1 gate2337( .a(N7272), .O(N8790) );
buf1 gate2338( .a(N7258), .O(N8793) );
buf1 gate2339( .a(N7258), .O(N8796) );
buf1 gate2340( .a(N7307), .O(N8799) );
buf1 gate2341( .a(N7288), .O(N8802) );
buf1 gate2342( .a(N7250), .O(N8805) );
buf1 gate2343( .a(N7272), .O(N8808) );
nand2 gate2344( .a(N8232), .b(N8233), .O(N8811) );
inv1 gate2345( .a(N7588), .O(N8814) );
inv1 gate2346( .a(N7591), .O(N8815) );
inv1 gate2347( .a(N7582), .O(N8816) );
inv1 gate2348( .a(N7585), .O(N8817) );
and2 gate2349( .a(N7620), .b(N3155), .O(N8818) );
and2 gate2350( .a(N3122), .b(N7609), .O(N8840) );
inv1 gate2351( .a(N7609), .O(N8857) );
and3 gate2352( .a(N6797), .b(N5740), .c(N8274), .O(N8861) );
and3 gate2353( .a(N5736), .b(N6800), .c(N8275), .O(N8862) );
and3 gate2354( .a(N6803), .b(N5751), .c(N8276), .O(N8863) );
and3 gate2355( .a(N5747), .b(N6806), .c(N8277), .O(N8864) );
and3 gate2356( .a(N6809), .b(N5762), .c(N8278), .O(N8865) );
and3 gate2357( .a(N5758), .b(N6812), .c(N8279), .O(N8866) );
inv1 gate2358( .a(N7655), .O(N8871) );
and2 gate2359( .a(N6833), .b(N7655), .O(N8874) );
and2 gate2360( .a(N7671), .b(N6867), .O(N8878) );
inv1 gate2361( .a(N8196), .O(N8879) );
nand2 gate2362( .a(N8196), .b(N8315), .O(N8880) );
inv1 gate2363( .a(N8200), .O(N8881) );
nand2 gate2364( .a(N8200), .b(N8317), .O(N8882) );
inv1 gate2365( .a(N8204), .O(N8883) );
nand2 gate2366( .a(N8204), .b(N8319), .O(N8884) );
inv1 gate2367( .a(N8208), .O(N8885) );
nand2 gate2368( .a(N8208), .b(N8321), .O(N8886) );
inv1 gate( .a(N3658),.O(N3658_NOT) );
inv1 gate( .a(N8323),.O(N8323_NOT));
and2 gate( .a(N3658_NOT), .b(p421), .O(EX1051) );
and2 gate( .a(N8323_NOT), .b(EX1051), .O(EX1052) );
and2 gate( .a(N3658), .b(p422), .O(EX1053) );
and2 gate( .a(N8323_NOT), .b(EX1053), .O(EX1054) );
and2 gate( .a(N3658_NOT), .b(p423), .O(EX1055) );
and2 gate( .a(N8323), .b(EX1055), .O(EX1056) );
and2 gate( .a(N3658), .b(p424), .O(EX1057) );
and2 gate( .a(N8323), .b(EX1057), .O(EX1058) );
or2  gate( .a(EX1052), .b(EX1054), .O(EX1059) );
or2  gate( .a(EX1056), .b(EX1059), .O(EX1060) );
or2  gate( .a(EX1058), .b(EX1060), .O(N8887) );
nand2 gate2370( .a(N4817), .b(N8325), .O(N8888) );
or4 gate2371( .a(N4544), .b(N8337), .c(N8338), .d(N8339), .O(N8898) );
or5 gate2372( .a(N4562), .b(N8348), .c(N8349), .d(N8350), .e(N8351), .O(N8902) );
or4 gate2373( .a(N4576), .b(N8369), .c(N8370), .d(N8371), .O(N8920) );
or2 gate2374( .a(N4581), .b(N8377), .O(N8924) );
or5 gate2375( .a(N4592), .b(N8378), .c(N8379), .d(N8380), .e(N8381), .O(N8927) );
or2 gate2376( .a(N4603), .b(N8392), .O(N8931) );
or2 gate2377( .a(N7825), .b(N8404), .O(N8943) );
or4 gate2378( .a(N4630), .b(N8409), .c(N8410), .d(N8411), .O(N8950) );
or5 gate2379( .a(N4637), .b(N8415), .c(N8416), .d(N8417), .e(N8418), .O(N8956) );
inv1 gate2380( .a(N7852), .O(N8959) );
and2 gate2381( .a(N3375), .b(N7852), .O(N8960) );
or4 gate2382( .a(N4656), .b(N8433), .c(N8434), .d(N8435), .O(N8963) );
or5 gate2383( .a(N4674), .b(N8447), .c(N8448), .d(N8449), .e(N8450), .O(N8966) );
and3 gate2384( .a(N7188), .b(N6083), .c(N8469), .O(N8991) );
and3 gate2385( .a(N6079), .b(N7191), .c(N8470), .O(N8992) );
or4 gate2386( .a(N4701), .b(N8488), .c(N8489), .d(N8490), .O(N8995) );
or2 gate2387( .a(N4706), .b(N8496), .O(N8996) );
or5 gate2388( .a(N4717), .b(N8500), .c(N8501), .d(N8502), .e(N8503), .O(N9001) );
or2 gate2389( .a(N4728), .b(N8516), .O(N9005) );
and3 gate2390( .a(N7334), .b(N6141), .c(N8537), .O(N9024) );
and3 gate2391( .a(N6137), .b(N7337), .c(N8538), .O(N9025) );
or4 gate2392( .a(N4756), .b(N8545), .c(N8546), .d(N8547), .O(N9029) );
or5 gate2393( .a(N4760), .b(N8551), .c(N8552), .d(N8553), .e(N8554), .O(N9035) );
and3 gate2394( .a(N7378), .b(N6170), .c(N8564), .O(N9053) );
and3 gate2395( .a(N6166), .b(N7381), .c(N8565), .O(N9054) );
nand2 gate2396( .a(N4303), .b(N8607), .O(N9064) );
nand2 gate2397( .a(N3507), .b(N8609), .O(N9065) );
inv1 gate2398( .a(N8114), .O(N9066) );
nand2 gate2399( .a(N8114), .b(N4795), .O(N9067) );
or2 gate2400( .a(N7613), .b(N6783), .O(N9068) );
inv1 gate2401( .a(N8117), .O(N9071) );
inv1 gate2402( .a(N8131), .O(N9072) );
nand2 gate2403( .a(N8131), .b(N6195), .O(N9073) );
inv1 gate2404( .a(N7613), .O(N9074) );
inv1 gate2405( .a(N8134), .O(N9077) );
or2 gate2406( .a(N7650), .b(N6865), .O(N9079) );
inv1 gate2407( .a(N8146), .O(N9082) );
inv1 gate2408( .a(N7650), .O(N9083) );
inv1 gate2409( .a(N8156), .O(N9086) );
inv1 gate2410( .a(N8166), .O(N9087) );
nand2 gate2411( .a(N8166), .b(N4813), .O(N9088) );
or2 gate2412( .a(N7659), .b(N6866), .O(N9089) );
inv1 gate2413( .a(N8169), .O(N9092) );
inv1 gate2414( .a(N8183), .O(N9093) );
inv1 gate( .a(N8183),.O(N8183_NOT) );
inv1 gate( .a(N6203),.O(N6203_NOT));
and2 gate( .a(N8183_NOT), .b(p425), .O(EX1061) );
and2 gate( .a(N6203_NOT), .b(EX1061), .O(EX1062) );
and2 gate( .a(N8183), .b(p426), .O(EX1063) );
and2 gate( .a(N6203_NOT), .b(EX1063), .O(EX1064) );
and2 gate( .a(N8183_NOT), .b(p427), .O(EX1065) );
and2 gate( .a(N6203), .b(EX1065), .O(EX1066) );
and2 gate( .a(N8183), .b(p428), .O(EX1067) );
and2 gate( .a(N6203), .b(EX1067), .O(EX1068) );
or2  gate( .a(EX1062), .b(EX1064), .O(EX1069) );
or2  gate( .a(EX1066), .b(EX1069), .O(EX1070) );
or2  gate( .a(EX1068), .b(EX1070), .O(N9094) );
inv1 gate2416( .a(N7659), .O(N9095) );
inv1 gate2417( .a(N8186), .O(N9098) );
or4 gate2418( .a(N4545), .b(N8340), .c(N8341), .d(N8342), .O(N9099) );
nor3 gate2419( .a(N4545), .b(N8343), .c(N8344), .O(N9103) );
or3 gate2420( .a(N4549), .b(N8345), .c(N8346), .O(N9107) );
nor2 gate2421( .a(N4549), .b(N8347), .O(N9111) );
or4 gate2422( .a(N4577), .b(N8372), .c(N8373), .d(N8374), .O(N9117) );
nor3 gate2423( .a(N4577), .b(N8375), .c(N8376), .O(N9127) );
nor3 gate2424( .a(N4597), .b(N8390), .c(N8391), .O(N9146) );
nor4 gate2425( .a(N4593), .b(N8385), .c(N8386), .d(N8387), .O(N9149) );
nand2 gate2426( .a(N7577), .b(N8733), .O(N9159) );
inv1 gate( .a(N7574),.O(N7574_NOT) );
inv1 gate( .a(N8734),.O(N8734_NOT));
and2 gate( .a(N7574_NOT), .b(p429), .O(EX1071) );
and2 gate( .a(N8734_NOT), .b(EX1071), .O(EX1072) );
and2 gate( .a(N7574), .b(p430), .O(EX1073) );
and2 gate( .a(N8734_NOT), .b(EX1073), .O(EX1074) );
and2 gate( .a(N7574_NOT), .b(p431), .O(EX1075) );
and2 gate( .a(N8734), .b(EX1075), .O(EX1076) );
and2 gate( .a(N7574), .b(p432), .O(EX1077) );
and2 gate( .a(N8734), .b(EX1077), .O(EX1078) );
or2  gate( .a(EX1072), .b(EX1074), .O(EX1079) );
or2  gate( .a(EX1076), .b(EX1079), .O(EX1080) );
or2  gate( .a(EX1078), .b(EX1080), .O(N9160) );
or4 gate2428( .a(N4657), .b(N8436), .c(N8437), .d(N8438), .O(N9161) );
nor3 gate2429( .a(N4657), .b(N8439), .c(N8440), .O(N9165) );
or3 gate2430( .a(N4661), .b(N8441), .c(N8442), .O(N9169) );
nor2 gate2431( .a(N4661), .b(N8443), .O(N9173) );
nand2 gate2432( .a(N7563), .b(N8753), .O(N9179) );
nand2 gate2433( .a(N7560), .b(N8754), .O(N9180) );
nand2 gate2434( .a(N7569), .b(N8755), .O(N9181) );
inv1 gate( .a(N7566),.O(N7566_NOT) );
inv1 gate( .a(N8756),.O(N8756_NOT));
and2 gate( .a(N7566_NOT), .b(p433), .O(EX1081) );
and2 gate( .a(N8756_NOT), .b(EX1081), .O(EX1082) );
and2 gate( .a(N7566), .b(p434), .O(EX1083) );
and2 gate( .a(N8756_NOT), .b(EX1083), .O(EX1084) );
and2 gate( .a(N7566_NOT), .b(p435), .O(EX1085) );
and2 gate( .a(N8756), .b(EX1085), .O(EX1086) );
and2 gate( .a(N7566), .b(p436), .O(EX1087) );
and2 gate( .a(N8756), .b(EX1087), .O(EX1088) );
or2  gate( .a(EX1082), .b(EX1084), .O(EX1089) );
or2  gate( .a(EX1086), .b(EX1089), .O(EX1090) );
or2  gate( .a(EX1088), .b(EX1090), .O(N9182) );
or4 gate2436( .a(N4702), .b(N8491), .c(N8492), .d(N8493), .O(N9183) );
nor3 gate2437( .a(N4702), .b(N8494), .c(N8495), .O(N9193) );
or4 gate2438( .a(N4722), .b(N8511), .c(N8512), .d(N8513), .O(N9203) );
or5 gate2439( .a(N4718), .b(N8504), .c(N8505), .d(N8506), .e(N8507), .O(N9206) );
nor3 gate2440( .a(N4722), .b(N8514), .c(N8515), .O(N9220) );
nor4 gate2441( .a(N4718), .b(N8508), .c(N8509), .d(N8510), .O(N9223) );
nand2 gate2442( .a(N7591), .b(N8814), .O(N9234) );
inv1 gate( .a(N7588),.O(N7588_NOT) );
inv1 gate( .a(N8815),.O(N8815_NOT));
and2 gate( .a(N7588_NOT), .b(p437), .O(EX1091) );
and2 gate( .a(N8815_NOT), .b(EX1091), .O(EX1092) );
and2 gate( .a(N7588), .b(p438), .O(EX1093) );
and2 gate( .a(N8815_NOT), .b(EX1093), .O(EX1094) );
and2 gate( .a(N7588_NOT), .b(p439), .O(EX1095) );
and2 gate( .a(N8815), .b(EX1095), .O(EX1096) );
and2 gate( .a(N7588), .b(p440), .O(EX1097) );
and2 gate( .a(N8815), .b(EX1097), .O(EX1098) );
or2  gate( .a(EX1092), .b(EX1094), .O(EX1099) );
or2  gate( .a(EX1096), .b(EX1099), .O(EX1100) );
or2  gate( .a(EX1098), .b(EX1100), .O(N9235) );
inv1 gate( .a(N7585),.O(N7585_NOT) );
inv1 gate( .a(N8816),.O(N8816_NOT));
and2 gate( .a(N7585_NOT), .b(p441), .O(EX1101) );
and2 gate( .a(N8816_NOT), .b(EX1101), .O(EX1102) );
and2 gate( .a(N7585), .b(p442), .O(EX1103) );
and2 gate( .a(N8816_NOT), .b(EX1103), .O(EX1104) );
and2 gate( .a(N7585_NOT), .b(p443), .O(EX1105) );
and2 gate( .a(N8816), .b(EX1105), .O(EX1106) );
and2 gate( .a(N7585), .b(p444), .O(EX1107) );
and2 gate( .a(N8816), .b(EX1107), .O(EX1108) );
or2  gate( .a(EX1102), .b(EX1104), .O(EX1109) );
or2  gate( .a(EX1106), .b(EX1109), .O(EX1110) );
or2  gate( .a(EX1108), .b(EX1110), .O(N9236) );
nand2 gate2445( .a(N7582), .b(N8817), .O(N9237) );
or2 gate2446( .a(N3159), .b(N8818), .O(N9238) );
or2 gate2447( .a(N3126), .b(N8840), .O(N9242) );
nand2 gate2448( .a(N8324), .b(N8888), .O(N9243) );
inv1 gate2449( .a(N8580), .O(N9244) );
inv1 gate2450( .a(N8583), .O(N9245) );
inv1 gate2451( .a(N8586), .O(N9246) );
inv1 gate2452( .a(N8589), .O(N9247) );
inv1 gate2453( .a(N8592), .O(N9248) );
inv1 gate2454( .a(N8595), .O(N9249) );
inv1 gate2455( .a(N8598), .O(N9250) );
inv1 gate2456( .a(N8601), .O(N9251) );
inv1 gate2457( .a(N8604), .O(N9252) );
nor2 gate2458( .a(N8861), .b(N8280), .O(N9256) );
nor2 gate2459( .a(N8862), .b(N8281), .O(N9257) );
nor2 gate2460( .a(N8863), .b(N8282), .O(N9258) );
inv1 gate( .a(N8864),.O(N8864_NOT) );
inv1 gate( .a(N8283),.O(N8283_NOT));
and2 gate( .a(N8864_NOT), .b(p445), .O(EX1111) );
and2 gate( .a(N8283_NOT), .b(EX1111), .O(EX1112) );
and2 gate( .a(N8864), .b(p446), .O(EX1113) );
and2 gate( .a(N8283_NOT), .b(EX1113), .O(EX1114) );
and2 gate( .a(N8864_NOT), .b(p447), .O(EX1115) );
and2 gate( .a(N8283), .b(EX1115), .O(EX1116) );
and2 gate( .a(N8864), .b(p448), .O(EX1117) );
and2 gate( .a(N8283), .b(EX1117), .O(EX1118) );
or2  gate( .a(EX1112), .b(EX1114), .O(EX1119) );
or2  gate( .a(EX1116), .b(EX1119), .O(EX1120) );
or2  gate( .a(EX1118), .b(EX1120), .O(N9259) );
nor2 gate2462( .a(N8865), .b(N8284), .O(N9260) );
nor2 gate2463( .a(N8866), .b(N8285), .O(N9261) );
inv1 gate2464( .a(N8627), .O(N9262) );
or2 gate2465( .a(N7649), .b(N8874), .O(N9265) );
or2 gate2466( .a(N7668), .b(N8878), .O(N9268) );
nand2 gate2467( .a(N7533), .b(N8879), .O(N9271) );
inv1 gate( .a(N7536),.O(N7536_NOT) );
inv1 gate( .a(N8881),.O(N8881_NOT));
and2 gate( .a(N7536_NOT), .b(p449), .O(EX1121) );
and2 gate( .a(N8881_NOT), .b(EX1121), .O(EX1122) );
and2 gate( .a(N7536), .b(p450), .O(EX1123) );
and2 gate( .a(N8881_NOT), .b(EX1123), .O(EX1124) );
and2 gate( .a(N7536_NOT), .b(p451), .O(EX1125) );
and2 gate( .a(N8881), .b(EX1125), .O(EX1126) );
and2 gate( .a(N7536), .b(p452), .O(EX1127) );
and2 gate( .a(N8881), .b(EX1127), .O(EX1128) );
or2  gate( .a(EX1122), .b(EX1124), .O(EX1129) );
or2  gate( .a(EX1126), .b(EX1129), .O(EX1130) );
or2  gate( .a(EX1128), .b(EX1130), .O(N9272) );
inv1 gate( .a(N7539),.O(N7539_NOT) );
inv1 gate( .a(N8883),.O(N8883_NOT));
and2 gate( .a(N7539_NOT), .b(p453), .O(EX1131) );
and2 gate( .a(N8883_NOT), .b(EX1131), .O(EX1132) );
and2 gate( .a(N7539), .b(p454), .O(EX1133) );
and2 gate( .a(N8883_NOT), .b(EX1133), .O(EX1134) );
and2 gate( .a(N7539_NOT), .b(p455), .O(EX1135) );
and2 gate( .a(N8883), .b(EX1135), .O(EX1136) );
and2 gate( .a(N7539), .b(p456), .O(EX1137) );
and2 gate( .a(N8883), .b(EX1137), .O(EX1138) );
or2  gate( .a(EX1132), .b(EX1134), .O(EX1139) );
or2  gate( .a(EX1136), .b(EX1139), .O(EX1140) );
or2  gate( .a(EX1138), .b(EX1140), .O(N9273) );
nand2 gate2470( .a(N7542), .b(N8885), .O(N9274) );
nand2 gate2471( .a(N8322), .b(N8887), .O(N9275) );
inv1 gate2472( .a(N8333), .O(N9276) );
and5 gate2473( .a(N6936), .b(N8326), .c(N6946), .d(N6929), .e(N6957), .O(N9280) );
and5 gate2474( .a(N367), .b(N8326), .c(N6946), .d(N6957), .e(N6936), .O(N9285) );
and4 gate2475( .a(N367), .b(N8326), .c(N6946), .d(N6957), .O(N9286) );
and3 gate2476( .a(N367), .b(N8326), .c(N6957), .O(N9287) );
and2 gate2477( .a(N367), .b(N8326), .O(N9288) );
inv1 gate2478( .a(N8660), .O(N9290) );
inv1 gate2479( .a(N8663), .O(N9292) );
inv1 gate2480( .a(N8666), .O(N9294) );
inv1 gate2481( .a(N8669), .O(N9296) );
inv1 gate( .a(N8672),.O(N8672_NOT) );
inv1 gate( .a(N5966),.O(N5966_NOT));
and2 gate( .a(N8672_NOT), .b(p457), .O(EX1141) );
and2 gate( .a(N5966_NOT), .b(EX1141), .O(EX1142) );
and2 gate( .a(N8672), .b(p458), .O(EX1143) );
and2 gate( .a(N5966_NOT), .b(EX1143), .O(EX1144) );
and2 gate( .a(N8672_NOT), .b(p459), .O(EX1145) );
and2 gate( .a(N5966), .b(EX1145), .O(EX1146) );
and2 gate( .a(N8672), .b(p460), .O(EX1147) );
and2 gate( .a(N5966), .b(EX1147), .O(EX1148) );
or2  gate( .a(EX1142), .b(EX1144), .O(EX1149) );
or2  gate( .a(EX1146), .b(EX1149), .O(EX1150) );
or2  gate( .a(EX1148), .b(EX1150), .O(N9297) );
inv1 gate2483( .a(N8672), .O(N9298) );
nand2 gate2484( .a(N8675), .b(N6969), .O(N9299) );
inv1 gate2485( .a(N8675), .O(N9300) );
inv1 gate2486( .a(N8365), .O(N9301) );
and5 gate2487( .a(N8358), .b(N7036), .c(N7020), .d(N7006), .e(N6998), .O(N9307) );
and4 gate2488( .a(N8358), .b(N7020), .c(N7006), .d(N7036), .O(N9314) );
and3 gate2489( .a(N8358), .b(N7020), .c(N7036), .O(N9315) );
and2 gate2490( .a(N8358), .b(N7036), .O(N9318) );
inv1 gate2491( .a(N8687), .O(N9319) );
inv1 gate2492( .a(N8699), .O(N9320) );
inv1 gate2493( .a(N8711), .O(N9321) );
inv1 gate2494( .a(N8714), .O(N9322) );
inv1 gate2495( .a(N8727), .O(N9323) );
inv1 gate2496( .a(N8730), .O(N9324) );
inv1 gate2497( .a(N8405), .O(N9326) );
and2 gate2498( .a(N8405), .b(N8412), .O(N9332) );
inv1 gate( .a(N4193),.O(N4193_NOT) );
inv1 gate( .a(N8960),.O(N8960_NOT));
and2 gate( .a(N4193_NOT), .b(p461), .O(EX1151) );
and2 gate( .a(N8960_NOT), .b(EX1151), .O(EX1152) );
and2 gate( .a(N4193), .b(p462), .O(EX1153) );
and2 gate( .a(N8960_NOT), .b(EX1153), .O(EX1154) );
and2 gate( .a(N4193_NOT), .b(p463), .O(EX1155) );
and2 gate( .a(N8960), .b(EX1155), .O(EX1156) );
and2 gate( .a(N4193), .b(p464), .O(EX1157) );
and2 gate( .a(N8960), .b(EX1157), .O(EX1158) );
or2  gate( .a(EX1152), .b(EX1154), .O(EX1159) );
or2  gate( .a(EX1156), .b(EX1159), .O(EX1160) );
or2  gate( .a(EX1158), .b(EX1160), .O(N9339) );
and2 gate2500( .a(N8430), .b(N8444), .O(N9344) );
inv1 gate2501( .a(N8735), .O(N9352) );
inv1 gate2502( .a(N8738), .O(N9354) );
inv1 gate2503( .a(N8741), .O(N9356) );
inv1 gate2504( .a(N8744), .O(N9358) );
nand2 gate2505( .a(N8747), .b(N6078), .O(N9359) );
inv1 gate2506( .a(N8747), .O(N9360) );
nand2 gate2507( .a(N8750), .b(N7187), .O(N9361) );
inv1 gate2508( .a(N8750), .O(N9362) );
inv1 gate2509( .a(N8471), .O(N9363) );
inv1 gate2510( .a(N8474), .O(N9364) );
inv1 gate2511( .a(N8477), .O(N9365) );
inv1 gate2512( .a(N8480), .O(N9366) );
inv1 gate( .a(N8991),.O(N8991_NOT) );
inv1 gate( .a(N8483),.O(N8483_NOT));
and2 gate( .a(N8991_NOT), .b(p465), .O(EX1161) );
and2 gate( .a(N8483_NOT), .b(EX1161), .O(EX1162) );
and2 gate( .a(N8991), .b(p466), .O(EX1163) );
and2 gate( .a(N8483_NOT), .b(EX1163), .O(EX1164) );
and2 gate( .a(N8991_NOT), .b(p467), .O(EX1165) );
and2 gate( .a(N8483), .b(EX1165), .O(EX1166) );
and2 gate( .a(N8991), .b(p468), .O(EX1167) );
and2 gate( .a(N8483), .b(EX1167), .O(EX1168) );
or2  gate( .a(EX1162), .b(EX1164), .O(EX1169) );
or2  gate( .a(EX1166), .b(EX1169), .O(EX1170) );
or2  gate( .a(EX1168), .b(EX1170), .O(N9367) );
nor2 gate2514( .a(N8992), .b(N8484), .O(N9368) );
and3 gate2515( .a(N7198), .b(N7194), .c(N8471), .O(N9369) );
and3 gate2516( .a(N8460), .b(N8457), .c(N8474), .O(N9370) );
and3 gate2517( .a(N7209), .b(N7205), .c(N8477), .O(N9371) );
and3 gate2518( .a(N8466), .b(N8463), .c(N8480), .O(N9372) );
inv1 gate2519( .a(N8497), .O(N9375) );
inv1 gate2520( .a(N8766), .O(N9381) );
inv1 gate2521( .a(N8778), .O(N9382) );
inv1 gate2522( .a(N8793), .O(N9383) );
inv1 gate2523( .a(N8796), .O(N9384) );
and2 gate2524( .a(N8485), .b(N8497), .O(N9385) );
inv1 gate2525( .a(N8525), .O(N9392) );
inv1 gate2526( .a(N8528), .O(N9393) );
inv1 gate2527( .a(N8531), .O(N9394) );
inv1 gate2528( .a(N8534), .O(N9395) );
and3 gate2529( .a(N7318), .b(N7314), .c(N8525), .O(N9396) );
and3 gate2530( .a(N8522), .b(N8519), .c(N8528), .O(N9397) );
and3 gate2531( .a(N6131), .b(N6127), .c(N8531), .O(N9398) );
and3 gate2532( .a(N7328), .b(N7325), .c(N8534), .O(N9399) );
inv1 gate( .a(N9024),.O(N9024_NOT) );
inv1 gate( .a(N8539),.O(N8539_NOT));
and2 gate( .a(N9024_NOT), .b(p469), .O(EX1171) );
and2 gate( .a(N8539_NOT), .b(EX1171), .O(EX1172) );
and2 gate( .a(N9024), .b(p470), .O(EX1173) );
and2 gate( .a(N8539_NOT), .b(EX1173), .O(EX1174) );
and2 gate( .a(N9024_NOT), .b(p471), .O(EX1175) );
and2 gate( .a(N8539), .b(EX1175), .O(EX1176) );
and2 gate( .a(N9024), .b(p472), .O(EX1177) );
and2 gate( .a(N8539), .b(EX1177), .O(EX1178) );
or2  gate( .a(EX1172), .b(EX1174), .O(EX1179) );
or2  gate( .a(EX1176), .b(EX1179), .O(EX1180) );
or2  gate( .a(EX1178), .b(EX1180), .O(N9400) );
nor2 gate2534( .a(N9025), .b(N8540), .O(N9401) );
inv1 gate2535( .a(N8541), .O(N9402) );
nand2 gate2536( .a(N8548), .b(N89), .O(N9407) );
and2 gate2537( .a(N8541), .b(N8548), .O(N9408) );
inv1 gate2538( .a(N8811), .O(N9412) );
inv1 gate2539( .a(N8566), .O(N9413) );
inv1 gate2540( .a(N8569), .O(N9414) );
inv1 gate2541( .a(N8572), .O(N9415) );
inv1 gate2542( .a(N8575), .O(N9416) );
inv1 gate( .a(N9053),.O(N9053_NOT) );
inv1 gate( .a(N8578),.O(N8578_NOT));
and2 gate( .a(N9053_NOT), .b(p473), .O(EX1181) );
and2 gate( .a(N8578_NOT), .b(EX1181), .O(EX1182) );
and2 gate( .a(N9053), .b(p474), .O(EX1183) );
and2 gate( .a(N8578_NOT), .b(EX1183), .O(EX1184) );
and2 gate( .a(N9053_NOT), .b(p475), .O(EX1185) );
and2 gate( .a(N8578), .b(EX1185), .O(EX1186) );
and2 gate( .a(N9053), .b(p476), .O(EX1187) );
and2 gate( .a(N8578), .b(EX1187), .O(EX1188) );
or2  gate( .a(EX1182), .b(EX1184), .O(EX1189) );
or2  gate( .a(EX1186), .b(EX1189), .O(EX1190) );
or2  gate( .a(EX1188), .b(EX1190), .O(N9417) );
nor2 gate2544( .a(N9054), .b(N8579), .O(N9418) );
and3 gate2545( .a(N7387), .b(N6177), .c(N8566), .O(N9419) );
and3 gate2546( .a(N8555), .b(N7384), .c(N8569), .O(N9420) );
and3 gate2547( .a(N7398), .b(N7394), .c(N8572), .O(N9421) );
and3 gate2548( .a(N8561), .b(N8558), .c(N8575), .O(N9422) );
buf1 gate2549( .a(N8326), .O(N9423) );
inv1 gate( .a(N9064),.O(N9064_NOT) );
inv1 gate( .a(N8608),.O(N8608_NOT));
and2 gate( .a(N9064_NOT), .b(p477), .O(EX1191) );
and2 gate( .a(N8608_NOT), .b(EX1191), .O(EX1192) );
and2 gate( .a(N9064), .b(p478), .O(EX1193) );
and2 gate( .a(N8608_NOT), .b(EX1193), .O(EX1194) );
and2 gate( .a(N9064_NOT), .b(p479), .O(EX1195) );
and2 gate( .a(N8608), .b(EX1195), .O(EX1196) );
and2 gate( .a(N9064), .b(p480), .O(EX1197) );
and2 gate( .a(N8608), .b(EX1197), .O(EX1198) );
or2  gate( .a(EX1192), .b(EX1194), .O(EX1199) );
or2  gate( .a(EX1196), .b(EX1199), .O(EX1200) );
or2  gate( .a(EX1198), .b(EX1200), .O(N9426) );
nand2 gate2551( .a(N9065), .b(N8610), .O(N9429) );
nand2 gate2552( .a(N3515), .b(N9066), .O(N9432) );
nand2 gate2553( .a(N4796), .b(N9072), .O(N9435) );
nand2 gate2554( .a(N3628), .b(N9087), .O(N9442) );
nand2 gate2555( .a(N4814), .b(N9093), .O(N9445) );
inv1 gate2556( .a(N8678), .O(N9454) );
inv1 gate2557( .a(N8681), .O(N9455) );
inv1 gate2558( .a(N8684), .O(N9456) );
inv1 gate2559( .a(N8690), .O(N9459) );
inv1 gate2560( .a(N8693), .O(N9460) );
inv1 gate2561( .a(N8696), .O(N9461) );
buf1 gate2562( .a(N8358), .O(N9462) );
inv1 gate2563( .a(N8702), .O(N9465) );
inv1 gate2564( .a(N8705), .O(N9466) );
inv1 gate2565( .a(N8708), .O(N9467) );
inv1 gate2566( .a(N8724), .O(N9468) );
buf1 gate2567( .a(N8358), .O(N9473) );
inv1 gate2568( .a(N8718), .O(N9476) );
inv1 gate2569( .a(N8721), .O(N9477) );
nand2 gate2570( .a(N9159), .b(N9160), .O(N9478) );
nand2 gate2571( .a(N9179), .b(N9180), .O(N9485) );
nand2 gate2572( .a(N9181), .b(N9182), .O(N9488) );
inv1 gate2573( .a(N8757), .O(N9493) );
inv1 gate2574( .a(N8760), .O(N9494) );
inv1 gate2575( .a(N8763), .O(N9495) );
inv1 gate2576( .a(N8769), .O(N9498) );
inv1 gate2577( .a(N8772), .O(N9499) );
inv1 gate2578( .a(N8775), .O(N9500) );
inv1 gate2579( .a(N8781), .O(N9505) );
inv1 gate2580( .a(N8784), .O(N9506) );
inv1 gate2581( .a(N8787), .O(N9507) );
inv1 gate2582( .a(N8790), .O(N9508) );
inv1 gate2583( .a(N8808), .O(N9509) );
inv1 gate2584( .a(N8799), .O(N9514) );
inv1 gate2585( .a(N8802), .O(N9515) );
inv1 gate2586( .a(N8805), .O(N9516) );
nand2 gate2587( .a(N9234), .b(N9235), .O(N9517) );
nand2 gate2588( .a(N9236), .b(N9237), .O(N9520) );
and2 gate2589( .a(N8943), .b(N8421), .O(N9526) );
and2 gate2590( .a(N8943), .b(N8421), .O(N9531) );
nand2 gate2591( .a(N9271), .b(N8880), .O(N9539) );
nand2 gate2592( .a(N9273), .b(N8884), .O(N9540) );
inv1 gate2593( .a(N9275), .O(N9541) );
and2 gate2594( .a(N8857), .b(N8254), .O(N9543) );
and2 gate2595( .a(N8871), .b(N8288), .O(N9551) );
nand2 gate2596( .a(N9272), .b(N8882), .O(N9555) );
nand2 gate2597( .a(N9274), .b(N8886), .O(N9556) );
inv1 gate2598( .a(N8898), .O(N9557) );
and2 gate2599( .a(N8902), .b(N8333), .O(N9560) );
inv1 gate2600( .a(N9099), .O(N9561) );
nand2 gate2601( .a(N9099), .b(N9290), .O(N9562) );
inv1 gate2602( .a(N9103), .O(N9563) );
nand2 gate2603( .a(N9103), .b(N9292), .O(N9564) );
inv1 gate2604( .a(N9107), .O(N9565) );
nand2 gate2605( .a(N9107), .b(N9294), .O(N9566) );
inv1 gate2606( .a(N9111), .O(N9567) );
nand2 gate2607( .a(N9111), .b(N9296), .O(N9568) );
nand2 gate2608( .a(N4844), .b(N9298), .O(N9569) );
nand2 gate2609( .a(N6207), .b(N9300), .O(N9570) );
inv1 gate2610( .a(N8920), .O(N9571) );
inv1 gate2611( .a(N8927), .O(N9575) );
and2 gate2612( .a(N8365), .b(N8927), .O(N9579) );
inv1 gate2613( .a(N8950), .O(N9581) );
inv1 gate2614( .a(N8956), .O(N9582) );
and2 gate2615( .a(N8405), .b(N8956), .O(N9585) );
and2 gate2616( .a(N8966), .b(N8430), .O(N9591) );
inv1 gate2617( .a(N9161), .O(N9592) );
nand2 gate2618( .a(N9161), .b(N9352), .O(N9593) );
inv1 gate2619( .a(N9165), .O(N9594) );
nand2 gate2620( .a(N9165), .b(N9354), .O(N9595) );
inv1 gate2621( .a(N9169), .O(N9596) );
inv1 gate( .a(N9169),.O(N9169_NOT) );
inv1 gate( .a(N9356),.O(N9356_NOT));
and2 gate( .a(N9169_NOT), .b(p481), .O(EX1201) );
and2 gate( .a(N9356_NOT), .b(EX1201), .O(EX1202) );
and2 gate( .a(N9169), .b(p482), .O(EX1203) );
and2 gate( .a(N9356_NOT), .b(EX1203), .O(EX1204) );
and2 gate( .a(N9169_NOT), .b(p483), .O(EX1205) );
and2 gate( .a(N9356), .b(EX1205), .O(EX1206) );
and2 gate( .a(N9169), .b(p484), .O(EX1207) );
and2 gate( .a(N9356), .b(EX1207), .O(EX1208) );
or2  gate( .a(EX1202), .b(EX1204), .O(EX1209) );
or2  gate( .a(EX1206), .b(EX1209), .O(EX1210) );
or2  gate( .a(EX1208), .b(EX1210), .O(N9597) );
inv1 gate2623( .a(N9173), .O(N9598) );
nand2 gate2624( .a(N9173), .b(N9358), .O(N9599) );
inv1 gate( .a(N4940),.O(N4940_NOT) );
inv1 gate( .a(N9360),.O(N9360_NOT));
and2 gate( .a(N4940_NOT), .b(p485), .O(EX1211) );
and2 gate( .a(N9360_NOT), .b(EX1211), .O(EX1212) );
and2 gate( .a(N4940), .b(p486), .O(EX1213) );
and2 gate( .a(N9360_NOT), .b(EX1213), .O(EX1214) );
and2 gate( .a(N4940_NOT), .b(p487), .O(EX1215) );
and2 gate( .a(N9360), .b(EX1215), .O(EX1216) );
and2 gate( .a(N4940), .b(p488), .O(EX1217) );
and2 gate( .a(N9360), .b(EX1217), .O(EX1218) );
or2  gate( .a(EX1212), .b(EX1214), .O(EX1219) );
or2  gate( .a(EX1216), .b(EX1219), .O(EX1220) );
or2  gate( .a(EX1218), .b(EX1220), .O(N9600) );
nand2 gate2626( .a(N6220), .b(N9362), .O(N9601) );
and3 gate2627( .a(N8457), .b(N7198), .c(N9363), .O(N9602) );
and3 gate2628( .a(N7194), .b(N8460), .c(N9364), .O(N9603) );
and3 gate2629( .a(N8463), .b(N7209), .c(N9365), .O(N9604) );
and3 gate2630( .a(N7205), .b(N8466), .c(N9366), .O(N9605) );
inv1 gate2631( .a(N9001), .O(N9608) );
and2 gate2632( .a(N8485), .b(N9001), .O(N9611) );
and3 gate2633( .a(N8519), .b(N7318), .c(N9392), .O(N9612) );
and3 gate2634( .a(N7314), .b(N8522), .c(N9393), .O(N9613) );
and3 gate2635( .a(N7325), .b(N6131), .c(N9394), .O(N9614) );
and3 gate2636( .a(N6127), .b(N7328), .c(N9395), .O(N9615) );
inv1 gate2637( .a(N9029), .O(N9616) );
inv1 gate2638( .a(N9035), .O(N9617) );
and2 gate2639( .a(N8541), .b(N9035), .O(N9618) );
and3 gate2640( .a(N7384), .b(N7387), .c(N9413), .O(N9621) );
and3 gate2641( .a(N6177), .b(N8555), .c(N9414), .O(N9622) );
and3 gate2642( .a(N8558), .b(N7398), .c(N9415), .O(N9623) );
and3 gate2643( .a(N7394), .b(N8561), .c(N9416), .O(N9624) );
or5 gate2644( .a(N4563), .b(N8352), .c(N8353), .d(N8354), .e(N9285), .O(N9626) );
or4 gate2645( .a(N4566), .b(N8355), .c(N8356), .d(N9286), .O(N9629) );
or3 gate2646( .a(N4570), .b(N8357), .c(N9287), .O(N9632) );
or2 gate2647( .a(N5960), .b(N9288), .O(N9635) );
nand2 gate2648( .a(N9067), .b(N9432), .O(N9642) );
inv1 gate2649( .a(N9068), .O(N9645) );
nand2 gate2650( .a(N9073), .b(N9435), .O(N9646) );
inv1 gate2651( .a(N9074), .O(N9649) );
nand2 gate2652( .a(N9257), .b(N9256), .O(N9650) );
nand2 gate2653( .a(N9259), .b(N9258), .O(N9653) );
nand2 gate2654( .a(N9261), .b(N9260), .O(N9656) );
inv1 gate2655( .a(N9079), .O(N9659) );
nand2 gate2656( .a(N9079), .b(N4809), .O(N9660) );
inv1 gate2657( .a(N9083), .O(N9661) );
nand2 gate2658( .a(N9083), .b(N6202), .O(N9662) );
nand2 gate2659( .a(N9088), .b(N9442), .O(N9663) );
inv1 gate2660( .a(N9089), .O(N9666) );
nand2 gate2661( .a(N9094), .b(N9445), .O(N9667) );
inv1 gate2662( .a(N9095), .O(N9670) );
or2 gate2663( .a(N8924), .b(N8393), .O(N9671) );
inv1 gate2664( .a(N9117), .O(N9674) );
inv1 gate2665( .a(N8924), .O(N9675) );
inv1 gate2666( .a(N9127), .O(N9678) );
or4 gate2667( .a(N4597), .b(N8388), .c(N8389), .d(N9315), .O(N9679) );
or2 gate2668( .a(N8931), .b(N9318), .O(N9682) );
or5 gate2669( .a(N4593), .b(N8382), .c(N8383), .d(N8384), .e(N9314), .O(N9685) );
inv1 gate2670( .a(N9146), .O(N9690) );
nand2 gate2671( .a(N9146), .b(N8717), .O(N9691) );
inv1 gate2672( .a(N8931), .O(N9692) );
inv1 gate2673( .a(N9149), .O(N9695) );
nand2 gate2674( .a(N9401), .b(N9400), .O(N9698) );
inv1 gate( .a(N9368),.O(N9368_NOT) );
inv1 gate( .a(N9367),.O(N9367_NOT));
and2 gate( .a(N9368_NOT), .b(p489), .O(EX1221) );
and2 gate( .a(N9367_NOT), .b(EX1221), .O(EX1222) );
and2 gate( .a(N9368), .b(p490), .O(EX1223) );
and2 gate( .a(N9367_NOT), .b(EX1223), .O(EX1224) );
and2 gate( .a(N9368_NOT), .b(p491), .O(EX1225) );
and2 gate( .a(N9367), .b(EX1225), .O(EX1226) );
and2 gate( .a(N9368), .b(p492), .O(EX1227) );
and2 gate( .a(N9367), .b(EX1227), .O(EX1228) );
or2  gate( .a(EX1222), .b(EX1224), .O(EX1229) );
or2  gate( .a(EX1226), .b(EX1229), .O(EX1230) );
or2  gate( .a(EX1228), .b(EX1230), .O(N9702) );
or2 gate2676( .a(N8996), .b(N8517), .O(N9707) );
inv1 gate2677( .a(N9183), .O(N9710) );
inv1 gate2678( .a(N8996), .O(N9711) );
inv1 gate2679( .a(N9193), .O(N9714) );
inv1 gate2680( .a(N9203), .O(N9715) );
nand2 gate2681( .a(N9203), .b(N6235), .O(N9716) );
or2 gate2682( .a(N9005), .b(N8518), .O(N9717) );
inv1 gate2683( .a(N9206), .O(N9720) );
inv1 gate2684( .a(N9220), .O(N9721) );
nand2 gate2685( .a(N9220), .b(N7573), .O(N9722) );
inv1 gate2686( .a(N9005), .O(N9723) );
inv1 gate2687( .a(N9223), .O(N9726) );
nand2 gate2688( .a(N9418), .b(N9417), .O(N9727) );
and2 gate2689( .a(N9268), .b(N8269), .O(N9732) );
nand2 gate2690( .a(N9581), .b(N9326), .O(N9733) );
and5 gate2691( .a(N89), .b(N9408), .c(N9332), .d(N8394), .e(N8421), .O(N9734) );
and5 gate2692( .a(N89), .b(N9408), .c(N9332), .d(N8394), .e(N8421), .O(N9735) );
and2 gate2693( .a(N9265), .b(N8262), .O(N9736) );
inv1 gate2694( .a(N9555), .O(N9737) );
inv1 gate2695( .a(N9556), .O(N9738) );
nand2 gate2696( .a(N9361), .b(N9601), .O(N9739) );
nand2 gate2697( .a(N9423), .b(N1115), .O(N9740) );
inv1 gate2698( .a(N9423), .O(N9741) );
nand2 gate2699( .a(N9299), .b(N9570), .O(N9742) );
and2 gate2700( .a(N8333), .b(N9280), .O(N9754) );
or2 gate2701( .a(N8898), .b(N9560), .O(N9758) );
nand2 gate2702( .a(N8660), .b(N9561), .O(N9762) );
nand2 gate2703( .a(N8663), .b(N9563), .O(N9763) );
nand2 gate2704( .a(N8666), .b(N9565), .O(N9764) );
nand2 gate2705( .a(N8669), .b(N9567), .O(N9765) );
nand2 gate2706( .a(N9297), .b(N9569), .O(N9766) );
and2 gate2707( .a(N9280), .b(N367), .O(N9767) );
nand2 gate2708( .a(N9557), .b(N9276), .O(N9768) );
inv1 gate2709( .a(N9307), .O(N9769) );
nand2 gate2710( .a(N9307), .b(N367), .O(N9773) );
inv1 gate( .a(N9571),.O(N9571_NOT) );
inv1 gate( .a(N9301),.O(N9301_NOT));
and2 gate( .a(N9571_NOT), .b(p493), .O(EX1231) );
and2 gate( .a(N9301_NOT), .b(EX1231), .O(EX1232) );
and2 gate( .a(N9571), .b(p494), .O(EX1233) );
and2 gate( .a(N9301_NOT), .b(EX1233), .O(EX1234) );
and2 gate( .a(N9571_NOT), .b(p495), .O(EX1235) );
and2 gate( .a(N9301), .b(EX1235), .O(EX1236) );
and2 gate( .a(N9571), .b(p496), .O(EX1237) );
and2 gate( .a(N9301), .b(EX1237), .O(EX1238) );
or2  gate( .a(EX1232), .b(EX1234), .O(EX1239) );
or2  gate( .a(EX1236), .b(EX1239), .O(EX1240) );
or2  gate( .a(EX1238), .b(EX1240), .O(N9774) );
and2 gate2712( .a(N8365), .b(N9307), .O(N9775) );
inv1 gate( .a(N8920),.O(N8920_NOT) );
inv1 gate( .a(N9579),.O(N9579_NOT));
and2 gate( .a(N8920_NOT), .b(p497), .O(EX1241) );
and2 gate( .a(N9579_NOT), .b(EX1241), .O(EX1242) );
and2 gate( .a(N8920), .b(p498), .O(EX1243) );
and2 gate( .a(N9579_NOT), .b(EX1243), .O(EX1244) );
and2 gate( .a(N8920_NOT), .b(p499), .O(EX1245) );
and2 gate( .a(N9579), .b(EX1245), .O(EX1246) );
and2 gate( .a(N8920), .b(p500), .O(EX1247) );
and2 gate( .a(N9579), .b(EX1247), .O(EX1248) );
or2  gate( .a(EX1242), .b(EX1244), .O(EX1249) );
or2  gate( .a(EX1246), .b(EX1249), .O(EX1250) );
or2  gate( .a(EX1248), .b(EX1250), .O(N9779) );
inv1 gate2714( .a(N9478), .O(N9784) );
inv1 gate( .a(N9616),.O(N9616_NOT) );
inv1 gate( .a(N9402),.O(N9402_NOT));
and2 gate( .a(N9616_NOT), .b(p501), .O(EX1251) );
and2 gate( .a(N9402_NOT), .b(EX1251), .O(EX1252) );
and2 gate( .a(N9616), .b(p502), .O(EX1253) );
and2 gate( .a(N9402_NOT), .b(EX1253), .O(EX1254) );
and2 gate( .a(N9616_NOT), .b(p503), .O(EX1255) );
and2 gate( .a(N9402), .b(EX1255), .O(EX1256) );
and2 gate( .a(N9616), .b(p504), .O(EX1257) );
and2 gate( .a(N9402), .b(EX1257), .O(EX1258) );
or2  gate( .a(EX1252), .b(EX1254), .O(EX1259) );
or2  gate( .a(EX1256), .b(EX1259), .O(EX1260) );
or2  gate( .a(EX1258), .b(EX1260), .O(N9785) );
inv1 gate( .a(N8950),.O(N8950_NOT) );
inv1 gate( .a(N9585),.O(N9585_NOT));
and2 gate( .a(N8950_NOT), .b(p505), .O(EX1261) );
and2 gate( .a(N9585_NOT), .b(EX1261), .O(EX1262) );
and2 gate( .a(N8950), .b(p506), .O(EX1263) );
and2 gate( .a(N9585_NOT), .b(EX1263), .O(EX1264) );
and2 gate( .a(N8950_NOT), .b(p507), .O(EX1265) );
and2 gate( .a(N9585), .b(EX1265), .O(EX1266) );
and2 gate( .a(N8950), .b(p508), .O(EX1267) );
and2 gate( .a(N9585), .b(EX1267), .O(EX1268) );
or2  gate( .a(EX1262), .b(EX1264), .O(EX1269) );
or2  gate( .a(EX1266), .b(EX1269), .O(EX1270) );
or2  gate( .a(EX1268), .b(EX1270), .O(N9786) );
and4 gate2717( .a(N89), .b(N9408), .c(N9332), .d(N8394), .O(N9790) );
inv1 gate( .a(N8963),.O(N8963_NOT) );
inv1 gate( .a(N9591),.O(N9591_NOT));
and2 gate( .a(N8963_NOT), .b(p509), .O(EX1271) );
and2 gate( .a(N9591_NOT), .b(EX1271), .O(EX1272) );
and2 gate( .a(N8963), .b(p510), .O(EX1273) );
and2 gate( .a(N9591_NOT), .b(EX1273), .O(EX1274) );
and2 gate( .a(N8963_NOT), .b(p511), .O(EX1275) );
and2 gate( .a(N9591), .b(EX1275), .O(EX1276) );
and2 gate( .a(N8963), .b(p512), .O(EX1277) );
and2 gate( .a(N9591), .b(EX1277), .O(EX1278) );
or2  gate( .a(EX1272), .b(EX1274), .O(EX1279) );
or2  gate( .a(EX1276), .b(EX1279), .O(EX1280) );
or2  gate( .a(EX1278), .b(EX1280), .O(N9791) );
inv1 gate( .a(N8735),.O(N8735_NOT) );
inv1 gate( .a(N9592),.O(N9592_NOT));
and2 gate( .a(N8735_NOT), .b(p513), .O(EX1281) );
and2 gate( .a(N9592_NOT), .b(EX1281), .O(EX1282) );
and2 gate( .a(N8735), .b(p514), .O(EX1283) );
and2 gate( .a(N9592_NOT), .b(EX1283), .O(EX1284) );
and2 gate( .a(N8735_NOT), .b(p515), .O(EX1285) );
and2 gate( .a(N9592), .b(EX1285), .O(EX1286) );
and2 gate( .a(N8735), .b(p516), .O(EX1287) );
and2 gate( .a(N9592), .b(EX1287), .O(EX1288) );
or2  gate( .a(EX1282), .b(EX1284), .O(EX1289) );
or2  gate( .a(EX1286), .b(EX1289), .O(EX1290) );
or2  gate( .a(EX1288), .b(EX1290), .O(N9795) );
nand2 gate2720( .a(N8738), .b(N9594), .O(N9796) );
nand2 gate2721( .a(N8741), .b(N9596), .O(N9797) );
nand2 gate2722( .a(N8744), .b(N9598), .O(N9798) );
nand2 gate2723( .a(N9359), .b(N9600), .O(N9799) );
nor2 gate2724( .a(N9602), .b(N9369), .O(N9800) );
nor2 gate2725( .a(N9603), .b(N9370), .O(N9801) );
nor2 gate2726( .a(N9604), .b(N9371), .O(N9802) );
nor2 gate2727( .a(N9605), .b(N9372), .O(N9803) );
inv1 gate2728( .a(N9485), .O(N9805) );
inv1 gate2729( .a(N9488), .O(N9806) );
or2 gate2730( .a(N8995), .b(N9611), .O(N9809) );
nor2 gate2731( .a(N9612), .b(N9396), .O(N9813) );
nor2 gate2732( .a(N9613), .b(N9397), .O(N9814) );
nor2 gate2733( .a(N9614), .b(N9398), .O(N9815) );
nor2 gate2734( .a(N9615), .b(N9399), .O(N9816) );
and2 gate2735( .a(N9617), .b(N9407), .O(N9817) );
inv1 gate( .a(N9029),.O(N9029_NOT) );
inv1 gate( .a(N9618),.O(N9618_NOT));
and2 gate( .a(N9029_NOT), .b(p517), .O(EX1291) );
and2 gate( .a(N9618_NOT), .b(EX1291), .O(EX1292) );
and2 gate( .a(N9029), .b(p518), .O(EX1293) );
and2 gate( .a(N9618_NOT), .b(EX1293), .O(EX1294) );
and2 gate( .a(N9029_NOT), .b(p519), .O(EX1295) );
and2 gate( .a(N9618), .b(EX1295), .O(EX1296) );
and2 gate( .a(N9029), .b(p520), .O(EX1297) );
and2 gate( .a(N9618), .b(EX1297), .O(EX1298) );
or2  gate( .a(EX1292), .b(EX1294), .O(EX1299) );
or2  gate( .a(EX1296), .b(EX1299), .O(EX1300) );
or2  gate( .a(EX1298), .b(EX1300), .O(N9820) );
inv1 gate2737( .a(N9517), .O(N9825) );
inv1 gate2738( .a(N9520), .O(N9826) );
nor2 gate2739( .a(N9621), .b(N9419), .O(N9827) );
nor2 gate2740( .a(N9622), .b(N9420), .O(N9828) );
inv1 gate( .a(N9623),.O(N9623_NOT) );
inv1 gate( .a(N9421),.O(N9421_NOT));
and2 gate( .a(N9623_NOT), .b(p521), .O(EX1301) );
and2 gate( .a(N9421_NOT), .b(EX1301), .O(EX1302) );
and2 gate( .a(N9623), .b(p522), .O(EX1303) );
and2 gate( .a(N9421_NOT), .b(EX1303), .O(EX1304) );
and2 gate( .a(N9623_NOT), .b(p523), .O(EX1305) );
and2 gate( .a(N9421), .b(EX1305), .O(EX1306) );
and2 gate( .a(N9623), .b(p524), .O(EX1307) );
and2 gate( .a(N9421), .b(EX1307), .O(EX1308) );
or2  gate( .a(EX1302), .b(EX1304), .O(EX1309) );
or2  gate( .a(EX1306), .b(EX1309), .O(EX1310) );
or2  gate( .a(EX1308), .b(EX1310), .O(N9829) );
nor2 gate2742( .a(N9624), .b(N9422), .O(N9830) );
inv1 gate2743( .a(N9426), .O(N9835) );
nand2 gate2744( .a(N9426), .b(N4789), .O(N9836) );
inv1 gate2745( .a(N9429), .O(N9837) );
nand2 gate2746( .a(N9429), .b(N4794), .O(N9838) );
nand2 gate2747( .a(N3625), .b(N9659), .O(N9846) );
nand2 gate2748( .a(N4810), .b(N9661), .O(N9847) );
inv1 gate2749( .a(N9462), .O(N9862) );
nand2 gate2750( .a(N7553), .b(N9690), .O(N9863) );
inv1 gate2751( .a(N9473), .O(N9866) );
inv1 gate( .a(N5030),.O(N5030_NOT) );
inv1 gate( .a(N9715),.O(N9715_NOT));
and2 gate( .a(N5030_NOT), .b(p525), .O(EX1311) );
and2 gate( .a(N9715_NOT), .b(EX1311), .O(EX1312) );
and2 gate( .a(N5030), .b(p526), .O(EX1313) );
and2 gate( .a(N9715_NOT), .b(EX1313), .O(EX1314) );
and2 gate( .a(N5030_NOT), .b(p527), .O(EX1315) );
and2 gate( .a(N9715), .b(EX1315), .O(EX1316) );
and2 gate( .a(N5030), .b(p528), .O(EX1317) );
and2 gate( .a(N9715), .b(EX1317), .O(EX1318) );
or2  gate( .a(EX1312), .b(EX1314), .O(EX1319) );
or2  gate( .a(EX1316), .b(EX1319), .O(EX1320) );
or2  gate( .a(EX1318), .b(EX1320), .O(N9873) );
nand2 gate2753( .a(N6236), .b(N9721), .O(N9876) );
nand2 gate2754( .a(N9795), .b(N9593), .O(N9890) );
nand2 gate2755( .a(N9797), .b(N9597), .O(N9891) );
inv1 gate2756( .a(N9799), .O(N9892) );
nand2 gate2757( .a(N871), .b(N9741), .O(N9893) );
nand2 gate2758( .a(N9762), .b(N9562), .O(N9894) );
inv1 gate( .a(N9764),.O(N9764_NOT) );
inv1 gate( .a(N9566),.O(N9566_NOT));
and2 gate( .a(N9764_NOT), .b(p529), .O(EX1321) );
and2 gate( .a(N9566_NOT), .b(EX1321), .O(EX1322) );
and2 gate( .a(N9764), .b(p530), .O(EX1323) );
and2 gate( .a(N9566_NOT), .b(EX1323), .O(EX1324) );
and2 gate( .a(N9764_NOT), .b(p531), .O(EX1325) );
and2 gate( .a(N9566), .b(EX1325), .O(EX1326) );
and2 gate( .a(N9764), .b(p532), .O(EX1327) );
and2 gate( .a(N9566), .b(EX1327), .O(EX1328) );
or2  gate( .a(EX1322), .b(EX1324), .O(EX1329) );
or2  gate( .a(EX1326), .b(EX1329), .O(EX1330) );
or2  gate( .a(EX1328), .b(EX1330), .O(N9895) );
inv1 gate2760( .a(N9766), .O(N9896) );
inv1 gate2761( .a(N9626), .O(N9897) );
nand2 gate2762( .a(N9626), .b(N9249), .O(N9898) );
inv1 gate2763( .a(N9629), .O(N9899) );
nand2 gate2764( .a(N9629), .b(N9250), .O(N9900) );
inv1 gate2765( .a(N9632), .O(N9901) );
nand2 gate2766( .a(N9632), .b(N9251), .O(N9902) );
inv1 gate2767( .a(N9635), .O(N9903) );
nand2 gate2768( .a(N9635), .b(N9252), .O(N9904) );
inv1 gate2769( .a(N9543), .O(N9905) );
inv1 gate2770( .a(N9650), .O(N9906) );
nand2 gate2771( .a(N9650), .b(N5769), .O(N9907) );
inv1 gate2772( .a(N9653), .O(N9908) );
nand2 gate2773( .a(N9653), .b(N5770), .O(N9909) );
inv1 gate2774( .a(N9656), .O(N9910) );
nand2 gate2775( .a(N9656), .b(N9262), .O(N9911) );
inv1 gate2776( .a(N9551), .O(N9917) );
nand2 gate2777( .a(N9763), .b(N9564), .O(N9923) );
inv1 gate( .a(N9765),.O(N9765_NOT) );
inv1 gate( .a(N9568),.O(N9568_NOT));
and2 gate( .a(N9765_NOT), .b(p533), .O(EX1331) );
and2 gate( .a(N9568_NOT), .b(EX1331), .O(EX1332) );
and2 gate( .a(N9765), .b(p534), .O(EX1333) );
and2 gate( .a(N9568_NOT), .b(EX1333), .O(EX1334) );
and2 gate( .a(N9765_NOT), .b(p535), .O(EX1335) );
and2 gate( .a(N9568), .b(EX1335), .O(EX1336) );
and2 gate( .a(N9765), .b(p536), .O(EX1337) );
and2 gate( .a(N9568), .b(EX1337), .O(EX1338) );
or2  gate( .a(EX1332), .b(EX1334), .O(EX1339) );
or2  gate( .a(EX1336), .b(EX1339), .O(EX1340) );
or2  gate( .a(EX1338), .b(EX1340), .O(N9924) );
or2 gate2779( .a(N8902), .b(N9767), .O(N9925) );
and2 gate2780( .a(N9575), .b(N9773), .O(N9932) );
and2 gate2781( .a(N9575), .b(N9769), .O(N9935) );
inv1 gate2782( .a(N9698), .O(N9938) );
nand2 gate2783( .a(N9698), .b(N9323), .O(N9939) );
nand2 gate2784( .a(N9796), .b(N9595), .O(N9945) );
nand2 gate2785( .a(N9798), .b(N9599), .O(N9946) );
inv1 gate2786( .a(N9702), .O(N9947) );
nand2 gate2787( .a(N9702), .b(N6102), .O(N9948) );
inv1 gate( .a(N9608),.O(N9608_NOT) );
inv1 gate( .a(N9375),.O(N9375_NOT));
and2 gate( .a(N9608_NOT), .b(p537), .O(EX1341) );
and2 gate( .a(N9375_NOT), .b(EX1341), .O(EX1342) );
and2 gate( .a(N9608), .b(p538), .O(EX1343) );
and2 gate( .a(N9375_NOT), .b(EX1343), .O(EX1344) );
and2 gate( .a(N9608_NOT), .b(p539), .O(EX1345) );
and2 gate( .a(N9375), .b(EX1345), .O(EX1346) );
and2 gate( .a(N9608), .b(p540), .O(EX1347) );
and2 gate( .a(N9375), .b(EX1347), .O(EX1348) );
or2  gate( .a(EX1342), .b(EX1344), .O(EX1349) );
or2  gate( .a(EX1346), .b(EX1349), .O(EX1350) );
or2  gate( .a(EX1348), .b(EX1350), .O(N9949) );
inv1 gate2789( .a(N9727), .O(N9953) );
nand2 gate2790( .a(N9727), .b(N9412), .O(N9954) );
nand2 gate2791( .a(N3502), .b(N9835), .O(N9955) );
nand2 gate2792( .a(N3510), .b(N9837), .O(N9956) );
inv1 gate2793( .a(N9642), .O(N9957) );
nand2 gate2794( .a(N9642), .b(N9645), .O(N9958) );
inv1 gate2795( .a(N9646), .O(N9959) );
nand2 gate2796( .a(N9646), .b(N9649), .O(N9960) );
nand2 gate2797( .a(N9660), .b(N9846), .O(N9961) );
nand2 gate2798( .a(N9662), .b(N9847), .O(N9964) );
inv1 gate2799( .a(N9663), .O(N9967) );
nand2 gate2800( .a(N9663), .b(N9666), .O(N9968) );
inv1 gate2801( .a(N9667), .O(N9969) );
nand2 gate2802( .a(N9667), .b(N9670), .O(N9970) );
inv1 gate2803( .a(N9671), .O(N9971) );
nand2 gate2804( .a(N9671), .b(N6213), .O(N9972) );
inv1 gate2805( .a(N9675), .O(N9973) );
nand2 gate2806( .a(N9675), .b(N7551), .O(N9974) );
inv1 gate2807( .a(N9679), .O(N9975) );
nand2 gate2808( .a(N9679), .b(N7552), .O(N9976) );
inv1 gate2809( .a(N9682), .O(N9977) );
inv1 gate2810( .a(N9685), .O(N9978) );
nand2 gate2811( .a(N9691), .b(N9863), .O(N9979) );
inv1 gate2812( .a(N9692), .O(N9982) );
nand2 gate2813( .a(N9814), .b(N9813), .O(N9983) );
nand2 gate2814( .a(N9816), .b(N9815), .O(N9986) );
nand2 gate2815( .a(N9801), .b(N9800), .O(N9989) );
nand2 gate2816( .a(N9803), .b(N9802), .O(N9992) );
inv1 gate2817( .a(N9707), .O(N9995) );
nand2 gate2818( .a(N9707), .b(N6231), .O(N9996) );
inv1 gate2819( .a(N9711), .O(N9997) );
nand2 gate2820( .a(N9711), .b(N7572), .O(N9998) );
nand2 gate2821( .a(N9716), .b(N9873), .O(N9999) );
inv1 gate2822( .a(N9717), .O(N10002) );
nand2 gate2823( .a(N9722), .b(N9876), .O(N10003) );
inv1 gate2824( .a(N9723), .O(N10006) );
nand2 gate2825( .a(N9830), .b(N9829), .O(N10007) );
nand2 gate2826( .a(N9828), .b(N9827), .O(N10010) );
and3 gate2827( .a(N9791), .b(N8307), .c(N8269), .O(N10013) );
and4 gate2828( .a(N9758), .b(N9344), .c(N8307), .d(N8269), .O(N10014) );
and5 gate2829( .a(N367), .b(N9754), .c(N9344), .d(N8307), .e(N8269), .O(N10015) );
and3 gate2830( .a(N9786), .b(N8394), .c(N8421), .O(N10016) );
and4 gate2831( .a(N9820), .b(N9332), .c(N8394), .d(N8421), .O(N10017) );
and3 gate2832( .a(N9786), .b(N8394), .c(N8421), .O(N10018) );
and4 gate2833( .a(N9820), .b(N9332), .c(N8394), .d(N8421), .O(N10019) );
and3 gate2834( .a(N9809), .b(N8298), .c(N8262), .O(N10020) );
and4 gate2835( .a(N9779), .b(N9385), .c(N8298), .d(N8262), .O(N10021) );
and5 gate2836( .a(N367), .b(N9775), .c(N9385), .d(N8298), .e(N8262), .O(N10022) );
inv1 gate2837( .a(N9945), .O(N10023) );
inv1 gate2838( .a(N9946), .O(N10024) );
nand2 gate2839( .a(N9740), .b(N9893), .O(N10025) );
inv1 gate2840( .a(N9923), .O(N10026) );
inv1 gate2841( .a(N9924), .O(N10028) );
nand2 gate2842( .a(N8595), .b(N9897), .O(N10032) );
inv1 gate( .a(N8598),.O(N8598_NOT) );
inv1 gate( .a(N9899),.O(N9899_NOT));
and2 gate( .a(N8598_NOT), .b(p541), .O(EX1351) );
and2 gate( .a(N9899_NOT), .b(EX1351), .O(EX1352) );
and2 gate( .a(N8598), .b(p542), .O(EX1353) );
and2 gate( .a(N9899_NOT), .b(EX1353), .O(EX1354) );
and2 gate( .a(N8598_NOT), .b(p543), .O(EX1355) );
and2 gate( .a(N9899), .b(EX1355), .O(EX1356) );
and2 gate( .a(N8598), .b(p544), .O(EX1357) );
and2 gate( .a(N9899), .b(EX1357), .O(EX1358) );
or2  gate( .a(EX1352), .b(EX1354), .O(EX1359) );
or2  gate( .a(EX1356), .b(EX1359), .O(EX1360) );
or2  gate( .a(EX1358), .b(EX1360), .O(N10033) );
nand2 gate2844( .a(N8601), .b(N9901), .O(N10034) );
nand2 gate2845( .a(N8604), .b(N9903), .O(N10035) );
nand2 gate2846( .a(N4803), .b(N9906), .O(N10036) );
nand2 gate2847( .a(N4806), .b(N9908), .O(N10037) );
nand2 gate2848( .a(N8627), .b(N9910), .O(N10038) );
and2 gate2849( .a(N9809), .b(N8298), .O(N10039) );
and3 gate2850( .a(N9779), .b(N9385), .c(N8298), .O(N10040) );
and4 gate2851( .a(N367), .b(N9775), .c(N9385), .d(N8298), .O(N10041) );
and2 gate2852( .a(N9779), .b(N9385), .O(N10042) );
and3 gate2853( .a(N367), .b(N9775), .c(N9385), .O(N10043) );
nand2 gate2854( .a(N8727), .b(N9938), .O(N10050) );
inv1 gate2855( .a(N9817), .O(N10053) );
inv1 gate( .a(N9817),.O(N9817_NOT) );
inv1 gate( .a(N9029),.O(N9029_NOT));
and2 gate( .a(N9817_NOT), .b(p545), .O(EX1361) );
and2 gate( .a(N9029_NOT), .b(EX1361), .O(EX1362) );
and2 gate( .a(N9817), .b(p546), .O(EX1363) );
and2 gate( .a(N9029_NOT), .b(EX1363), .O(EX1364) );
and2 gate( .a(N9817_NOT), .b(p547), .O(EX1365) );
and2 gate( .a(N9029), .b(EX1365), .O(EX1366) );
and2 gate( .a(N9817), .b(p548), .O(EX1367) );
and2 gate( .a(N9029), .b(EX1367), .O(EX1368) );
or2  gate( .a(EX1362), .b(EX1364), .O(EX1369) );
or2  gate( .a(EX1366), .b(EX1369), .O(EX1370) );
or2  gate( .a(EX1368), .b(EX1370), .O(N10054) );
and2 gate2857( .a(N9786), .b(N8394), .O(N10055) );
and3 gate2858( .a(N9820), .b(N9332), .c(N8394), .O(N10056) );
and2 gate2859( .a(N9791), .b(N8307), .O(N10057) );
and3 gate2860( .a(N9758), .b(N9344), .c(N8307), .O(N10058) );
and4 gate2861( .a(N367), .b(N9754), .c(N9344), .d(N8307), .O(N10059) );
and2 gate2862( .a(N9758), .b(N9344), .O(N10060) );
and3 gate2863( .a(N367), .b(N9754), .c(N9344), .O(N10061) );
nand2 gate2864( .a(N4997), .b(N9947), .O(N10062) );
nand2 gate2865( .a(N8811), .b(N9953), .O(N10067) );
nand2 gate2866( .a(N9955), .b(N9836), .O(N10070) );
nand2 gate2867( .a(N9956), .b(N9838), .O(N10073) );
nand2 gate2868( .a(N9068), .b(N9957), .O(N10076) );
nand2 gate2869( .a(N9074), .b(N9959), .O(N10077) );
nand2 gate2870( .a(N9089), .b(N9967), .O(N10082) );
nand2 gate2871( .a(N9095), .b(N9969), .O(N10083) );
inv1 gate( .a(N4871),.O(N4871_NOT) );
inv1 gate( .a(N9971),.O(N9971_NOT));
and2 gate( .a(N4871_NOT), .b(p549), .O(EX1371) );
and2 gate( .a(N9971_NOT), .b(EX1371), .O(EX1372) );
and2 gate( .a(N4871), .b(p550), .O(EX1373) );
and2 gate( .a(N9971_NOT), .b(EX1373), .O(EX1374) );
and2 gate( .a(N4871_NOT), .b(p551), .O(EX1375) );
and2 gate( .a(N9971), .b(EX1375), .O(EX1376) );
and2 gate( .a(N4871), .b(p552), .O(EX1377) );
and2 gate( .a(N9971), .b(EX1377), .O(EX1378) );
or2  gate( .a(EX1372), .b(EX1374), .O(EX1379) );
or2  gate( .a(EX1376), .b(EX1379), .O(EX1380) );
or2  gate( .a(EX1378), .b(EX1380), .O(N10084) );
nand2 gate2873( .a(N6214), .b(N9973), .O(N10085) );
nand2 gate2874( .a(N6217), .b(N9975), .O(N10086) );
nand2 gate2875( .a(N5027), .b(N9995), .O(N10093) );
nand2 gate2876( .a(N6232), .b(N9997), .O(N10094) );
or5 gate2877( .a(N9238), .b(N9732), .c(N10013), .d(N10014), .e(N10015), .O(N10101) );
or5 gate2878( .a(N9339), .b(N9526), .c(N10016), .d(N10017), .e(N9734), .O(N10102) );
or5 gate2879( .a(N9339), .b(N9531), .c(N10018), .d(N10019), .e(N9735), .O(N10103) );
or5 gate2880( .a(N9242), .b(N9736), .c(N10020), .d(N10021), .e(N10022), .O(N10104) );
and2 gate2881( .a(N9925), .b(N9894), .O(N10105) );
inv1 gate( .a(N9925),.O(N9925_NOT) );
inv1 gate( .a(N9895),.O(N9895_NOT));
and2 gate( .a(N9925_NOT), .b(p553), .O(EX1381) );
and2 gate( .a(N9895_NOT), .b(EX1381), .O(EX1382) );
and2 gate( .a(N9925), .b(p554), .O(EX1383) );
and2 gate( .a(N9895_NOT), .b(EX1383), .O(EX1384) );
and2 gate( .a(N9925_NOT), .b(p555), .O(EX1385) );
and2 gate( .a(N9895), .b(EX1385), .O(EX1386) );
and2 gate( .a(N9925), .b(p556), .O(EX1387) );
and2 gate( .a(N9895), .b(EX1387), .O(EX1388) );
or2  gate( .a(EX1382), .b(EX1384), .O(EX1389) );
or2  gate( .a(EX1386), .b(EX1389), .O(EX1390) );
or2  gate( .a(EX1388), .b(EX1390), .O(N10106) );
inv1 gate( .a(N9925),.O(N9925_NOT) );
inv1 gate( .a(N9896),.O(N9896_NOT));
and2 gate( .a(N9925_NOT), .b(p557), .O(EX1391) );
and2 gate( .a(N9896_NOT), .b(EX1391), .O(EX1392) );
and2 gate( .a(N9925), .b(p558), .O(EX1393) );
and2 gate( .a(N9896_NOT), .b(EX1393), .O(EX1394) );
and2 gate( .a(N9925_NOT), .b(p559), .O(EX1395) );
and2 gate( .a(N9896), .b(EX1395), .O(EX1396) );
and2 gate( .a(N9925), .b(p560), .O(EX1397) );
and2 gate( .a(N9896), .b(EX1397), .O(EX1398) );
or2  gate( .a(EX1392), .b(EX1394), .O(EX1399) );
or2  gate( .a(EX1396), .b(EX1399), .O(EX1400) );
or2  gate( .a(EX1398), .b(EX1400), .O(N10107) );
and2 gate2884( .a(N9925), .b(N8253), .O(N10108) );
nand2 gate2885( .a(N10032), .b(N9898), .O(N10109) );
nand2 gate2886( .a(N10033), .b(N9900), .O(N10110) );
nand2 gate2887( .a(N10034), .b(N9902), .O(N10111) );
nand2 gate2888( .a(N10035), .b(N9904), .O(N10112) );
nand2 gate2889( .a(N10036), .b(N9907), .O(N10113) );
nand2 gate2890( .a(N10037), .b(N9909), .O(N10114) );
nand2 gate2891( .a(N10038), .b(N9911), .O(N10115) );
or4 gate2892( .a(N9265), .b(N10039), .c(N10040), .d(N10041), .O(N10116) );
or3 gate2893( .a(N9809), .b(N10042), .c(N10043), .O(N10119) );
inv1 gate2894( .a(N9925), .O(N10124) );
and2 gate2895( .a(N9768), .b(N9925), .O(N10130) );
inv1 gate2896( .a(N9932), .O(N10131) );
inv1 gate2897( .a(N9935), .O(N10132) );
and2 gate2898( .a(N9932), .b(N8920), .O(N10133) );
nand2 gate2899( .a(N10050), .b(N9939), .O(N10134) );
inv1 gate2900( .a(N9983), .O(N10135) );
nand2 gate2901( .a(N9983), .b(N9324), .O(N10136) );
inv1 gate2902( .a(N9986), .O(N10137) );
nand2 gate2903( .a(N9986), .b(N9784), .O(N10138) );
and2 gate2904( .a(N9785), .b(N10053), .O(N10139) );
or4 gate2905( .a(N8943), .b(N10055), .c(N10056), .d(N9790), .O(N10140) );
or4 gate2906( .a(N9268), .b(N10057), .c(N10058), .d(N10059), .O(N10141) );
or3 gate2907( .a(N9791), .b(N10060), .c(N10061), .O(N10148) );
nand2 gate2908( .a(N10062), .b(N9948), .O(N10155) );
inv1 gate2909( .a(N9989), .O(N10156) );
nand2 gate2910( .a(N9989), .b(N9805), .O(N10157) );
inv1 gate2911( .a(N9992), .O(N10158) );
nand2 gate2912( .a(N9992), .b(N9806), .O(N10159) );
inv1 gate2913( .a(N9949), .O(N10160) );
nand2 gate2914( .a(N10067), .b(N9954), .O(N10161) );
inv1 gate2915( .a(N10007), .O(N10162) );
nand2 gate2916( .a(N10007), .b(N9825), .O(N10163) );
inv1 gate2917( .a(N10010), .O(N10164) );
nand2 gate2918( .a(N10010), .b(N9826), .O(N10165) );
nand2 gate2919( .a(N10076), .b(N9958), .O(N10170) );
nand2 gate2920( .a(N10077), .b(N9960), .O(N10173) );
inv1 gate2921( .a(N9961), .O(N10176) );
nand2 gate2922( .a(N9961), .b(N9082), .O(N10177) );
inv1 gate2923( .a(N9964), .O(N10178) );
nand2 gate2924( .a(N9964), .b(N9086), .O(N10179) );
inv1 gate( .a(N10082),.O(N10082_NOT) );
inv1 gate( .a(N9968),.O(N9968_NOT));
and2 gate( .a(N10082_NOT), .b(p561), .O(EX1401) );
and2 gate( .a(N9968_NOT), .b(EX1401), .O(EX1402) );
and2 gate( .a(N10082), .b(p562), .O(EX1403) );
and2 gate( .a(N9968_NOT), .b(EX1403), .O(EX1404) );
and2 gate( .a(N10082_NOT), .b(p563), .O(EX1405) );
and2 gate( .a(N9968), .b(EX1405), .O(EX1406) );
and2 gate( .a(N10082), .b(p564), .O(EX1407) );
and2 gate( .a(N9968), .b(EX1407), .O(EX1408) );
or2  gate( .a(EX1402), .b(EX1404), .O(EX1409) );
or2  gate( .a(EX1406), .b(EX1409), .O(EX1410) );
or2  gate( .a(EX1408), .b(EX1410), .O(N10180) );
nand2 gate2926( .a(N10083), .b(N9970), .O(N10183) );
nand2 gate2927( .a(N9972), .b(N10084), .O(N10186) );
nand2 gate2928( .a(N9974), .b(N10085), .O(N10189) );
nand2 gate2929( .a(N9976), .b(N10086), .O(N10192) );
inv1 gate2930( .a(N9979), .O(N10195) );
nand2 gate2931( .a(N9979), .b(N9982), .O(N10196) );
nand2 gate2932( .a(N9996), .b(N10093), .O(N10197) );
nand2 gate2933( .a(N9998), .b(N10094), .O(N10200) );
inv1 gate2934( .a(N9999), .O(N10203) );
nand2 gate2935( .a(N9999), .b(N10002), .O(N10204) );
inv1 gate2936( .a(N10003), .O(N10205) );
nand2 gate2937( .a(N10003), .b(N10006), .O(N10206) );
nand2 gate2938( .a(N10070), .b(N4308), .O(N10212) );
nand2 gate2939( .a(N10073), .b(N4313), .O(N10213) );
and2 gate2940( .a(N9774), .b(N10131), .O(N10230) );
nand2 gate2941( .a(N8730), .b(N10135), .O(N10231) );
inv1 gate( .a(N9478),.O(N9478_NOT) );
inv1 gate( .a(N10137),.O(N10137_NOT));
and2 gate( .a(N9478_NOT), .b(p565), .O(EX1411) );
and2 gate( .a(N10137_NOT), .b(EX1411), .O(EX1412) );
and2 gate( .a(N9478), .b(p566), .O(EX1413) );
and2 gate( .a(N10137_NOT), .b(EX1413), .O(EX1414) );
and2 gate( .a(N9478_NOT), .b(p567), .O(EX1415) );
and2 gate( .a(N10137), .b(EX1415), .O(EX1416) );
and2 gate( .a(N9478), .b(p568), .O(EX1417) );
and2 gate( .a(N10137), .b(EX1417), .O(EX1418) );
or2  gate( .a(EX1412), .b(EX1414), .O(EX1419) );
or2  gate( .a(EX1416), .b(EX1419), .O(EX1420) );
or2  gate( .a(EX1418), .b(EX1420), .O(N10232) );
or2 gate2943( .a(N10139), .b(N10054), .O(N10233) );
inv1 gate( .a(N7100),.O(N7100_NOT) );
inv1 gate( .a(N10140),.O(N10140_NOT));
and2 gate( .a(N7100_NOT), .b(p569), .O(EX1421) );
and2 gate( .a(N10140_NOT), .b(EX1421), .O(EX1422) );
and2 gate( .a(N7100), .b(p570), .O(EX1423) );
and2 gate( .a(N10140_NOT), .b(EX1423), .O(EX1424) );
and2 gate( .a(N7100_NOT), .b(p571), .O(EX1425) );
and2 gate( .a(N10140), .b(EX1425), .O(EX1426) );
and2 gate( .a(N7100), .b(p572), .O(EX1427) );
and2 gate( .a(N10140), .b(EX1427), .O(EX1428) );
or2  gate( .a(EX1422), .b(EX1424), .O(EX1429) );
or2  gate( .a(EX1426), .b(EX1429), .O(EX1430) );
or2  gate( .a(EX1428), .b(EX1430), .O(N10234) );
nand2 gate2945( .a(N9485), .b(N10156), .O(N10237) );
nand2 gate2946( .a(N9488), .b(N10158), .O(N10238) );
nand2 gate2947( .a(N9517), .b(N10162), .O(N10239) );
nand2 gate2948( .a(N9520), .b(N10164), .O(N10240) );
inv1 gate2949( .a(N10070), .O(N10241) );
inv1 gate2950( .a(N10073), .O(N10242) );
nand2 gate2951( .a(N8146), .b(N10176), .O(N10247) );
nand2 gate2952( .a(N8156), .b(N10178), .O(N10248) );
nand2 gate2953( .a(N9692), .b(N10195), .O(N10259) );
nand2 gate2954( .a(N9717), .b(N10203), .O(N10264) );
nand2 gate2955( .a(N9723), .b(N10205), .O(N10265) );
and2 gate2956( .a(N10026), .b(N10124), .O(N10266) );
and2 gate2957( .a(N10028), .b(N10124), .O(N10267) );
and2 gate2958( .a(N9742), .b(N10124), .O(N10268) );
and2 gate2959( .a(N6923), .b(N10124), .O(N10269) );
nand2 gate2960( .a(N6762), .b(N10116), .O(N10270) );
inv1 gate( .a(N3061),.O(N3061_NOT) );
inv1 gate( .a(N10241),.O(N10241_NOT));
and2 gate( .a(N3061_NOT), .b(p573), .O(EX1431) );
and2 gate( .a(N10241_NOT), .b(EX1431), .O(EX1432) );
and2 gate( .a(N3061), .b(p574), .O(EX1433) );
and2 gate( .a(N10241_NOT), .b(EX1433), .O(EX1434) );
and2 gate( .a(N3061_NOT), .b(p575), .O(EX1435) );
and2 gate( .a(N10241), .b(EX1435), .O(EX1436) );
and2 gate( .a(N3061), .b(p576), .O(EX1437) );
and2 gate( .a(N10241), .b(EX1437), .O(EX1438) );
or2  gate( .a(EX1432), .b(EX1434), .O(EX1439) );
or2  gate( .a(EX1436), .b(EX1439), .O(EX1440) );
or2  gate( .a(EX1438), .b(EX1440), .O(N10271) );
nand2 gate2962( .a(N3064), .b(N10242), .O(N10272) );
buf1 gate2963( .a(N10116), .O(N10273) );
and5 gate2964( .a(N10141), .b(N5728), .c(N5707), .d(N5718), .e(N5697), .O(N10278) );
and4 gate2965( .a(N10141), .b(N5728), .c(N5707), .d(N5718), .O(N10279) );
and3 gate2966( .a(N10141), .b(N5728), .c(N5718), .O(N10280) );
and2 gate2967( .a(N10141), .b(N5728), .O(N10281) );
and2 gate2968( .a(N6784), .b(N10141), .O(N10282) );
inv1 gate2969( .a(N10119), .O(N10283) );
and5 gate2970( .a(N10148), .b(N5936), .c(N5915), .d(N5926), .e(N5905), .O(N10287) );
and4 gate2971( .a(N10148), .b(N5936), .c(N5915), .d(N5926), .O(N10288) );
and3 gate2972( .a(N10148), .b(N5936), .c(N5926), .O(N10289) );
and2 gate2973( .a(N10148), .b(N5936), .O(N10290) );
and2 gate2974( .a(N6881), .b(N10148), .O(N10291) );
and2 gate2975( .a(N8898), .b(N10124), .O(N10292) );
nand2 gate2976( .a(N10231), .b(N10136), .O(N10293) );
nand2 gate2977( .a(N10232), .b(N10138), .O(N10294) );
nand2 gate2978( .a(N8412), .b(N10233), .O(N10295) );
and2 gate2979( .a(N8959), .b(N10234), .O(N10296) );
nand2 gate2980( .a(N10237), .b(N10157), .O(N10299) );
nand2 gate2981( .a(N10238), .b(N10159), .O(N10300) );
or2 gate2982( .a(N10230), .b(N10133), .O(N10301) );
nand2 gate2983( .a(N10239), .b(N10163), .O(N10306) );
nand2 gate2984( .a(N10240), .b(N10165), .O(N10307) );
buf1 gate2985( .a(N10148), .O(N10308) );
buf1 gate2986( .a(N10141), .O(N10311) );
inv1 gate2987( .a(N10170), .O(N10314) );
nand2 gate2988( .a(N10170), .b(N9071), .O(N10315) );
inv1 gate2989( .a(N10173), .O(N10316) );
nand2 gate2990( .a(N10173), .b(N9077), .O(N10317) );
nand2 gate2991( .a(N10247), .b(N10177), .O(N10318) );
nand2 gate2992( .a(N10248), .b(N10179), .O(N10321) );
inv1 gate2993( .a(N10180), .O(N10324) );
nand2 gate2994( .a(N10180), .b(N9092), .O(N10325) );
inv1 gate2995( .a(N10183), .O(N10326) );
nand2 gate2996( .a(N10183), .b(N9098), .O(N10327) );
inv1 gate2997( .a(N10186), .O(N10328) );
nand2 gate2998( .a(N10186), .b(N9674), .O(N10329) );
inv1 gate2999( .a(N10189), .O(N10330) );
nand2 gate3000( .a(N10189), .b(N9678), .O(N10331) );
inv1 gate3001( .a(N10192), .O(N10332) );
nand2 gate3002( .a(N10192), .b(N9977), .O(N10333) );
nand2 gate3003( .a(N10259), .b(N10196), .O(N10334) );
inv1 gate3004( .a(N10197), .O(N10337) );
nand2 gate3005( .a(N10197), .b(N9710), .O(N10338) );
inv1 gate3006( .a(N10200), .O(N10339) );
nand2 gate3007( .a(N10200), .b(N9714), .O(N10340) );
nand2 gate3008( .a(N10264), .b(N10204), .O(N10341) );
nand2 gate3009( .a(N10265), .b(N10206), .O(N10344) );
or2 gate3010( .a(N10266), .b(N10105), .O(N10350) );
or2 gate3011( .a(N10267), .b(N10106), .O(N10351) );
or2 gate3012( .a(N10268), .b(N10107), .O(N10352) );
or2 gate3013( .a(N10269), .b(N10108), .O(N10353) );
and2 gate3014( .a(N8857), .b(N10270), .O(N10354) );
nand2 gate3015( .a(N10271), .b(N10212), .O(N10357) );
nand2 gate3016( .a(N10272), .b(N10213), .O(N10360) );
inv1 gate( .a(N7620),.O(N7620_NOT) );
inv1 gate( .a(N10282),.O(N10282_NOT));
and2 gate( .a(N7620_NOT), .b(p577), .O(EX1441) );
and2 gate( .a(N10282_NOT), .b(EX1441), .O(EX1442) );
and2 gate( .a(N7620), .b(p578), .O(EX1443) );
and2 gate( .a(N10282_NOT), .b(EX1443), .O(EX1444) );
and2 gate( .a(N7620_NOT), .b(p579), .O(EX1445) );
and2 gate( .a(N10282), .b(EX1445), .O(EX1446) );
and2 gate( .a(N7620), .b(p580), .O(EX1447) );
and2 gate( .a(N10282), .b(EX1447), .O(EX1448) );
or2  gate( .a(EX1442), .b(EX1444), .O(EX1449) );
or2  gate( .a(EX1446), .b(EX1449), .O(EX1450) );
or2  gate( .a(EX1448), .b(EX1450), .O(N10367) );
or2 gate3018( .a(N7671), .b(N10291), .O(N10375) );
or2 gate3019( .a(N10292), .b(N10130), .O(N10381) );
and4 gate3020( .a(N10114), .b(N10134), .c(N10293), .d(N10294), .O(N10388) );
and2 gate3021( .a(N9582), .b(N10295), .O(N10391) );
and4 gate3022( .a(N10113), .b(N10115), .c(N10299), .d(N10300), .O(N10399) );
and4 gate3023( .a(N10155), .b(N10161), .c(N10306), .d(N10307), .O(N10402) );
or5 gate3024( .a(N3229), .b(N6888), .c(N6889), .d(N6890), .e(N10287), .O(N10406) );
or4 gate3025( .a(N3232), .b(N6891), .c(N6892), .d(N10288), .O(N10409) );
or3 gate3026( .a(N3236), .b(N6893), .c(N10289), .O(N10412) );
inv1 gate( .a(N3241),.O(N3241_NOT) );
inv1 gate( .a(N10290),.O(N10290_NOT));
and2 gate( .a(N3241_NOT), .b(p581), .O(EX1451) );
and2 gate( .a(N10290_NOT), .b(EX1451), .O(EX1452) );
and2 gate( .a(N3241), .b(p582), .O(EX1453) );
and2 gate( .a(N10290_NOT), .b(EX1453), .O(EX1454) );
and2 gate( .a(N3241_NOT), .b(p583), .O(EX1455) );
and2 gate( .a(N10290), .b(EX1455), .O(EX1456) );
and2 gate( .a(N3241), .b(p584), .O(EX1457) );
and2 gate( .a(N10290), .b(EX1457), .O(EX1458) );
or2  gate( .a(EX1452), .b(EX1454), .O(EX1459) );
or2  gate( .a(EX1456), .b(EX1459), .O(EX1460) );
or2  gate( .a(EX1458), .b(EX1460), .O(N10415) );
or5 gate3028( .a(N3137), .b(N6791), .c(N6792), .d(N6793), .e(N10278), .O(N10419) );
or4 gate3029( .a(N3140), .b(N6794), .c(N6795), .d(N10279), .O(N10422) );
or3 gate3030( .a(N3144), .b(N6796), .c(N10280), .O(N10425) );
or2 gate3031( .a(N3149), .b(N10281), .O(N10428) );
nand2 gate3032( .a(N8117), .b(N10314), .O(N10431) );
nand2 gate3033( .a(N8134), .b(N10316), .O(N10432) );
nand2 gate3034( .a(N8169), .b(N10324), .O(N10437) );
nand2 gate3035( .a(N8186), .b(N10326), .O(N10438) );
nand2 gate3036( .a(N9117), .b(N10328), .O(N10439) );
nand2 gate3037( .a(N9127), .b(N10330), .O(N10440) );
inv1 gate( .a(N9682),.O(N9682_NOT) );
inv1 gate( .a(N10332),.O(N10332_NOT));
and2 gate( .a(N9682_NOT), .b(p585), .O(EX1461) );
and2 gate( .a(N10332_NOT), .b(EX1461), .O(EX1462) );
and2 gate( .a(N9682), .b(p586), .O(EX1463) );
and2 gate( .a(N10332_NOT), .b(EX1463), .O(EX1464) );
and2 gate( .a(N9682_NOT), .b(p587), .O(EX1465) );
and2 gate( .a(N10332), .b(EX1465), .O(EX1466) );
and2 gate( .a(N9682), .b(p588), .O(EX1467) );
and2 gate( .a(N10332), .b(EX1467), .O(EX1468) );
or2  gate( .a(EX1462), .b(EX1464), .O(EX1469) );
or2  gate( .a(EX1466), .b(EX1469), .O(EX1470) );
or2  gate( .a(EX1468), .b(EX1470), .O(N10441) );
nand2 gate3039( .a(N9183), .b(N10337), .O(N10444) );
nand2 gate3040( .a(N9193), .b(N10339), .O(N10445) );
inv1 gate3041( .a(N10296), .O(N10450) );
inv1 gate( .a(N10296),.O(N10296_NOT) );
inv1 gate( .a(N4193),.O(N4193_NOT));
and2 gate( .a(N10296_NOT), .b(p589), .O(EX1471) );
and2 gate( .a(N4193_NOT), .b(EX1471), .O(EX1472) );
and2 gate( .a(N10296), .b(p590), .O(EX1473) );
and2 gate( .a(N4193_NOT), .b(EX1473), .O(EX1474) );
and2 gate( .a(N10296_NOT), .b(p591), .O(EX1475) );
and2 gate( .a(N4193), .b(EX1475), .O(EX1476) );
and2 gate( .a(N10296), .b(p592), .O(EX1477) );
and2 gate( .a(N4193), .b(EX1477), .O(EX1478) );
or2  gate( .a(EX1472), .b(EX1474), .O(EX1479) );
or2  gate( .a(EX1476), .b(EX1479), .O(EX1480) );
or2  gate( .a(EX1478), .b(EX1480), .O(N10451) );
inv1 gate3043( .a(N10308), .O(N10455) );
nand2 gate3044( .a(N10308), .b(N8242), .O(N10456) );
inv1 gate3045( .a(N10311), .O(N10465) );
nand2 gate3046( .a(N10311), .b(N8247), .O(N10466) );
inv1 gate3047( .a(N10273), .O(N10479) );
inv1 gate3048( .a(N10301), .O(N10497) );
nand2 gate3049( .a(N10431), .b(N10315), .O(N10509) );
nand2 gate3050( .a(N10432), .b(N10317), .O(N10512) );
inv1 gate3051( .a(N10318), .O(N10515) );
nand2 gate3052( .a(N10318), .b(N8632), .O(N10516) );
inv1 gate3053( .a(N10321), .O(N10517) );
nand2 gate3054( .a(N10321), .b(N8637), .O(N10518) );
nand2 gate3055( .a(N10437), .b(N10325), .O(N10519) );
nand2 gate3056( .a(N10438), .b(N10327), .O(N10522) );
inv1 gate( .a(N10439),.O(N10439_NOT) );
inv1 gate( .a(N10329),.O(N10329_NOT));
and2 gate( .a(N10439_NOT), .b(p593), .O(EX1481) );
and2 gate( .a(N10329_NOT), .b(EX1481), .O(EX1482) );
and2 gate( .a(N10439), .b(p594), .O(EX1483) );
and2 gate( .a(N10329_NOT), .b(EX1483), .O(EX1484) );
and2 gate( .a(N10439_NOT), .b(p595), .O(EX1485) );
and2 gate( .a(N10329), .b(EX1485), .O(EX1486) );
and2 gate( .a(N10439), .b(p596), .O(EX1487) );
and2 gate( .a(N10329), .b(EX1487), .O(EX1488) );
or2  gate( .a(EX1482), .b(EX1484), .O(EX1489) );
or2  gate( .a(EX1486), .b(EX1489), .O(EX1490) );
or2  gate( .a(EX1488), .b(EX1490), .O(N10525) );
nand2 gate3058( .a(N10440), .b(N10331), .O(N10528) );
nand2 gate3059( .a(N10441), .b(N10333), .O(N10531) );
inv1 gate3060( .a(N10334), .O(N10534) );
nand2 gate3061( .a(N10334), .b(N9695), .O(N10535) );
nand2 gate3062( .a(N10444), .b(N10338), .O(N10536) );
nand2 gate3063( .a(N10445), .b(N10340), .O(N10539) );
inv1 gate3064( .a(N10341), .O(N10542) );
nand2 gate3065( .a(N10341), .b(N9720), .O(N10543) );
inv1 gate3066( .a(N10344), .O(N10544) );
nand2 gate3067( .a(N10344), .b(N9726), .O(N10545) );
and2 gate3068( .a(N5631), .b(N10450), .O(N10546) );
inv1 gate3069( .a(N10391), .O(N10547) );
inv1 gate( .a(N10391),.O(N10391_NOT) );
inv1 gate( .a(N8950),.O(N8950_NOT));
and2 gate( .a(N10391_NOT), .b(p597), .O(EX1491) );
and2 gate( .a(N8950_NOT), .b(EX1491), .O(EX1492) );
and2 gate( .a(N10391), .b(p598), .O(EX1493) );
and2 gate( .a(N8950_NOT), .b(EX1493), .O(EX1494) );
and2 gate( .a(N10391_NOT), .b(p599), .O(EX1495) );
and2 gate( .a(N8950), .b(EX1495), .O(EX1496) );
and2 gate( .a(N10391), .b(p600), .O(EX1497) );
and2 gate( .a(N8950), .b(EX1497), .O(EX1498) );
or2  gate( .a(EX1492), .b(EX1494), .O(EX1499) );
or2  gate( .a(EX1496), .b(EX1499), .O(EX1500) );
or2  gate( .a(EX1498), .b(EX1500), .O(N10548) );
inv1 gate( .a(N5165),.O(N5165_NOT) );
inv1 gate( .a(N10367),.O(N10367_NOT));
and2 gate( .a(N5165_NOT), .b(p601), .O(EX1501) );
and2 gate( .a(N10367_NOT), .b(EX1501), .O(EX1502) );
and2 gate( .a(N5165), .b(p602), .O(EX1503) );
and2 gate( .a(N10367_NOT), .b(EX1503), .O(EX1504) );
and2 gate( .a(N5165_NOT), .b(p603), .O(EX1505) );
and2 gate( .a(N10367), .b(EX1505), .O(EX1506) );
and2 gate( .a(N5165), .b(p604), .O(EX1507) );
and2 gate( .a(N10367), .b(EX1507), .O(EX1508) );
or2  gate( .a(EX1502), .b(EX1504), .O(EX1509) );
or2  gate( .a(EX1506), .b(EX1509), .O(EX1510) );
or2  gate( .a(EX1508), .b(EX1510), .O(N10549) );
inv1 gate3072( .a(N10354), .O(N10550) );
and2 gate3073( .a(N10354), .b(N3126), .O(N10551) );
nand2 gate3074( .a(N7411), .b(N10455), .O(N10552) );
and2 gate3075( .a(N10375), .b(N9539), .O(N10553) );
and2 gate3076( .a(N10375), .b(N9540), .O(N10554) );
and2 gate3077( .a(N10375), .b(N9541), .O(N10555) );
and2 gate3078( .a(N10375), .b(N6761), .O(N10556) );
inv1 gate3079( .a(N10406), .O(N10557) );
nand2 gate3080( .a(N10406), .b(N8243), .O(N10558) );
inv1 gate3081( .a(N10409), .O(N10559) );
nand2 gate3082( .a(N10409), .b(N8244), .O(N10560) );
inv1 gate3083( .a(N10412), .O(N10561) );
nand2 gate3084( .a(N10412), .b(N8245), .O(N10562) );
inv1 gate3085( .a(N10415), .O(N10563) );
nand2 gate3086( .a(N10415), .b(N8246), .O(N10564) );
nand2 gate3087( .a(N7426), .b(N10465), .O(N10565) );
inv1 gate3088( .a(N10419), .O(N10566) );
nand2 gate3089( .a(N10419), .b(N8248), .O(N10567) );
inv1 gate3090( .a(N10422), .O(N10568) );
nand2 gate3091( .a(N10422), .b(N8249), .O(N10569) );
inv1 gate3092( .a(N10425), .O(N10570) );
nand2 gate3093( .a(N10425), .b(N8250), .O(N10571) );
inv1 gate3094( .a(N10428), .O(N10572) );
nand2 gate3095( .a(N10428), .b(N8251), .O(N10573) );
inv1 gate3096( .a(N10399), .O(N10574) );
inv1 gate3097( .a(N10402), .O(N10575) );
inv1 gate3098( .a(N10388), .O(N10576) );
and3 gate3099( .a(N10399), .b(N10402), .c(N10388), .O(N10577) );
and3 gate3100( .a(N10360), .b(N9543), .c(N10273), .O(N10581) );
and3 gate3101( .a(N10357), .b(N9905), .c(N10273), .O(N10582) );
inv1 gate3102( .a(N10367), .O(N10583) );
and2 gate3103( .a(N10367), .b(N5735), .O(N10587) );
inv1 gate( .a(N10367),.O(N10367_NOT) );
inv1 gate( .a(N3135),.O(N3135_NOT));
and2 gate( .a(N10367_NOT), .b(p605), .O(EX1511) );
and2 gate( .a(N3135_NOT), .b(EX1511), .O(EX1512) );
and2 gate( .a(N10367), .b(p606), .O(EX1513) );
and2 gate( .a(N3135_NOT), .b(EX1513), .O(EX1514) );
and2 gate( .a(N10367_NOT), .b(p607), .O(EX1515) );
and2 gate( .a(N3135), .b(EX1515), .O(EX1516) );
and2 gate( .a(N10367), .b(p608), .O(EX1517) );
and2 gate( .a(N3135), .b(EX1517), .O(EX1518) );
or2  gate( .a(EX1512), .b(EX1514), .O(EX1519) );
or2  gate( .a(EX1516), .b(EX1519), .O(EX1520) );
or2  gate( .a(EX1518), .b(EX1520), .O(N10588) );
inv1 gate3105( .a(N10375), .O(N10589) );
and5 gate3106( .a(N10381), .b(N7180), .c(N7159), .d(N7170), .e(N7149), .O(N10594) );
and4 gate3107( .a(N10381), .b(N7180), .c(N7159), .d(N7170), .O(N10595) );
and3 gate3108( .a(N10381), .b(N7180), .c(N7170), .O(N10596) );
inv1 gate( .a(N10381),.O(N10381_NOT) );
inv1 gate( .a(N7180),.O(N7180_NOT));
and2 gate( .a(N10381_NOT), .b(p609), .O(EX1521) );
and2 gate( .a(N7180_NOT), .b(EX1521), .O(EX1522) );
and2 gate( .a(N10381), .b(p610), .O(EX1523) );
and2 gate( .a(N7180_NOT), .b(EX1523), .O(EX1524) );
and2 gate( .a(N10381_NOT), .b(p611), .O(EX1525) );
and2 gate( .a(N7180), .b(EX1525), .O(EX1526) );
and2 gate( .a(N10381), .b(p612), .O(EX1527) );
and2 gate( .a(N7180), .b(EX1527), .O(EX1528) );
or2  gate( .a(EX1522), .b(EX1524), .O(EX1529) );
or2  gate( .a(EX1526), .b(EX1529), .O(EX1530) );
or2  gate( .a(EX1528), .b(EX1530), .O(N10597) );
and2 gate3110( .a(N8444), .b(N10381), .O(N10598) );
buf1 gate3111( .a(N10381), .O(N10602) );
nand2 gate3112( .a(N7479), .b(N10515), .O(N10609) );
nand2 gate3113( .a(N7491), .b(N10517), .O(N10610) );
inv1 gate( .a(N9149),.O(N9149_NOT) );
inv1 gate( .a(N10534),.O(N10534_NOT));
and2 gate( .a(N9149_NOT), .b(p613), .O(EX1531) );
and2 gate( .a(N10534_NOT), .b(EX1531), .O(EX1532) );
and2 gate( .a(N9149), .b(p614), .O(EX1533) );
and2 gate( .a(N10534_NOT), .b(EX1533), .O(EX1534) );
and2 gate( .a(N9149_NOT), .b(p615), .O(EX1535) );
and2 gate( .a(N10534), .b(EX1535), .O(EX1536) );
and2 gate( .a(N9149), .b(p616), .O(EX1537) );
and2 gate( .a(N10534), .b(EX1537), .O(EX1538) );
or2  gate( .a(EX1532), .b(EX1534), .O(EX1539) );
or2  gate( .a(EX1536), .b(EX1539), .O(EX1540) );
or2  gate( .a(EX1538), .b(EX1540), .O(N10621) );
nand2 gate3115( .a(N9206), .b(N10542), .O(N10626) );
nand2 gate3116( .a(N9223), .b(N10544), .O(N10627) );
or2 gate3117( .a(N10546), .b(N10451), .O(N10628) );
inv1 gate( .a(N9733),.O(N9733_NOT) );
inv1 gate( .a(N10547),.O(N10547_NOT));
and2 gate( .a(N9733_NOT), .b(p617), .O(EX1541) );
and2 gate( .a(N10547_NOT), .b(EX1541), .O(EX1542) );
and2 gate( .a(N9733), .b(p618), .O(EX1543) );
and2 gate( .a(N10547_NOT), .b(EX1543), .O(EX1544) );
and2 gate( .a(N9733_NOT), .b(p619), .O(EX1545) );
and2 gate( .a(N10547), .b(EX1545), .O(EX1546) );
and2 gate( .a(N9733), .b(p620), .O(EX1547) );
and2 gate( .a(N10547), .b(EX1547), .O(EX1548) );
or2  gate( .a(EX1542), .b(EX1544), .O(EX1549) );
or2  gate( .a(EX1546), .b(EX1549), .O(EX1550) );
or2  gate( .a(EX1548), .b(EX1550), .O(N10629) );
inv1 gate( .a(N5166),.O(N5166_NOT) );
inv1 gate( .a(N10550),.O(N10550_NOT));
and2 gate( .a(N5166_NOT), .b(p621), .O(EX1551) );
and2 gate( .a(N10550_NOT), .b(EX1551), .O(EX1552) );
and2 gate( .a(N5166), .b(p622), .O(EX1553) );
and2 gate( .a(N10550_NOT), .b(EX1553), .O(EX1554) );
and2 gate( .a(N5166_NOT), .b(p623), .O(EX1555) );
and2 gate( .a(N10550), .b(EX1555), .O(EX1556) );
and2 gate( .a(N5166), .b(p624), .O(EX1557) );
and2 gate( .a(N10550), .b(EX1557), .O(EX1558) );
or2  gate( .a(EX1552), .b(EX1554), .O(EX1559) );
or2  gate( .a(EX1556), .b(EX1559), .O(EX1560) );
or2  gate( .a(EX1558), .b(EX1560), .O(N10631) );
nand2 gate3120( .a(N10552), .b(N10456), .O(N10632) );
nand2 gate3121( .a(N7414), .b(N10557), .O(N10637) );
nand2 gate3122( .a(N7417), .b(N10559), .O(N10638) );
nand2 gate3123( .a(N7420), .b(N10561), .O(N10639) );
nand2 gate3124( .a(N7423), .b(N10563), .O(N10640) );
nand2 gate3125( .a(N10565), .b(N10466), .O(N10641) );
nand2 gate3126( .a(N7429), .b(N10566), .O(N10642) );
nand2 gate3127( .a(N7432), .b(N10568), .O(N10643) );
nand2 gate3128( .a(N7435), .b(N10570), .O(N10644) );
nand2 gate3129( .a(N7438), .b(N10572), .O(N10645) );
and3 gate3130( .a(N886), .b(N887), .c(N10577), .O(N10647) );
and3 gate3131( .a(N10360), .b(N8857), .c(N10479), .O(N10648) );
and3 gate3132( .a(N10357), .b(N7609), .c(N10479), .O(N10649) );
or2 gate3133( .a(N8966), .b(N10598), .O(N10652) );
or5 gate3134( .a(N4675), .b(N8451), .c(N8452), .d(N8453), .e(N10594), .O(N10659) );
or4 gate3135( .a(N4678), .b(N8454), .c(N8455), .d(N10595), .O(N10662) );
or3 gate3136( .a(N4682), .b(N8456), .c(N10596), .O(N10665) );
or2 gate3137( .a(N4687), .b(N10597), .O(N10668) );
inv1 gate3138( .a(N10509), .O(N10671) );
nand2 gate3139( .a(N10509), .b(N8615), .O(N10672) );
inv1 gate3140( .a(N10512), .O(N10673) );
nand2 gate3141( .a(N10512), .b(N8624), .O(N10674) );
nand2 gate3142( .a(N10609), .b(N10516), .O(N10675) );
nand2 gate3143( .a(N10610), .b(N10518), .O(N10678) );
inv1 gate3144( .a(N10519), .O(N10681) );
nand2 gate3145( .a(N10519), .b(N8644), .O(N10682) );
inv1 gate3146( .a(N10522), .O(N10683) );
nand2 gate3147( .a(N10522), .b(N8653), .O(N10684) );
inv1 gate3148( .a(N10525), .O(N10685) );
nand2 gate3149( .a(N10525), .b(N9454), .O(N10686) );
inv1 gate3150( .a(N10528), .O(N10687) );
nand2 gate3151( .a(N10528), .b(N9459), .O(N10688) );
inv1 gate3152( .a(N10531), .O(N10689) );
nand2 gate3153( .a(N10531), .b(N9978), .O(N10690) );
nand2 gate3154( .a(N10621), .b(N10535), .O(N10691) );
inv1 gate3155( .a(N10536), .O(N10694) );
nand2 gate3156( .a(N10536), .b(N9493), .O(N10695) );
inv1 gate3157( .a(N10539), .O(N10696) );
nand2 gate3158( .a(N10539), .b(N9498), .O(N10697) );
nand2 gate3159( .a(N10626), .b(N10543), .O(N10698) );
nand2 gate3160( .a(N10627), .b(N10545), .O(N10701) );
or2 gate3161( .a(N10629), .b(N10548), .O(N10704) );
inv1 gate( .a(N3159),.O(N3159_NOT) );
inv1 gate( .a(N10583),.O(N10583_NOT));
and2 gate( .a(N3159_NOT), .b(p625), .O(EX1561) );
and2 gate( .a(N10583_NOT), .b(EX1561), .O(EX1562) );
and2 gate( .a(N3159), .b(p626), .O(EX1563) );
and2 gate( .a(N10583_NOT), .b(EX1563), .O(EX1564) );
and2 gate( .a(N3159_NOT), .b(p627), .O(EX1565) );
and2 gate( .a(N10583), .b(EX1565), .O(EX1566) );
and2 gate( .a(N3159), .b(p628), .O(EX1567) );
and2 gate( .a(N10583), .b(EX1567), .O(EX1568) );
or2  gate( .a(EX1562), .b(EX1564), .O(EX1569) );
or2  gate( .a(EX1566), .b(EX1569), .O(EX1570) );
or2  gate( .a(EX1568), .b(EX1570), .O(N10705) );
or2 gate3163( .a(N10631), .b(N10551), .O(N10706) );
and2 gate3164( .a(N9737), .b(N10589), .O(N10707) );
and2 gate3165( .a(N9738), .b(N10589), .O(N10708) );
and2 gate3166( .a(N9243), .b(N10589), .O(N10709) );
and2 gate3167( .a(N5892), .b(N10589), .O(N10710) );
nand2 gate3168( .a(N10637), .b(N10558), .O(N10711) );
nand2 gate3169( .a(N10638), .b(N10560), .O(N10712) );
nand2 gate3170( .a(N10639), .b(N10562), .O(N10713) );
inv1 gate( .a(N10640),.O(N10640_NOT) );
inv1 gate( .a(N10564),.O(N10564_NOT));
and2 gate( .a(N10640_NOT), .b(p629), .O(EX1571) );
and2 gate( .a(N10564_NOT), .b(EX1571), .O(EX1572) );
and2 gate( .a(N10640), .b(p630), .O(EX1573) );
and2 gate( .a(N10564_NOT), .b(EX1573), .O(EX1574) );
and2 gate( .a(N10640_NOT), .b(p631), .O(EX1575) );
and2 gate( .a(N10564), .b(EX1575), .O(EX1576) );
and2 gate( .a(N10640), .b(p632), .O(EX1577) );
and2 gate( .a(N10564), .b(EX1577), .O(EX1578) );
or2  gate( .a(EX1572), .b(EX1574), .O(EX1579) );
or2  gate( .a(EX1576), .b(EX1579), .O(EX1580) );
or2  gate( .a(EX1578), .b(EX1580), .O(N10714) );
nand2 gate3172( .a(N10642), .b(N10567), .O(N10715) );
nand2 gate3173( .a(N10643), .b(N10569), .O(N10716) );
nand2 gate3174( .a(N10644), .b(N10571), .O(N10717) );
inv1 gate( .a(N10645),.O(N10645_NOT) );
inv1 gate( .a(N10573),.O(N10573_NOT));
and2 gate( .a(N10645_NOT), .b(p633), .O(EX1581) );
and2 gate( .a(N10573_NOT), .b(EX1581), .O(EX1582) );
and2 gate( .a(N10645), .b(p634), .O(EX1583) );
and2 gate( .a(N10573_NOT), .b(EX1583), .O(EX1584) );
and2 gate( .a(N10645_NOT), .b(p635), .O(EX1585) );
and2 gate( .a(N10573), .b(EX1585), .O(EX1586) );
and2 gate( .a(N10645), .b(p636), .O(EX1587) );
and2 gate( .a(N10573), .b(EX1587), .O(EX1588) );
or2  gate( .a(EX1582), .b(EX1584), .O(EX1589) );
or2  gate( .a(EX1586), .b(EX1589), .O(EX1590) );
or2  gate( .a(EX1588), .b(EX1590), .O(N10718) );
inv1 gate3176( .a(N10602), .O(N10719) );
nand2 gate3177( .a(N10602), .b(N9244), .O(N10720) );
inv1 gate3178( .a(N10647), .O(N10729) );
and2 gate3179( .a(N5178), .b(N10583), .O(N10730) );
and2 gate3180( .a(N2533), .b(N10583), .O(N10731) );
nand2 gate3181( .a(N7447), .b(N10671), .O(N10737) );
nand2 gate3182( .a(N7465), .b(N10673), .O(N10738) );
or4 gate3183( .a(N10648), .b(N10649), .c(N10581), .d(N10582), .O(N10739) );
nand2 gate3184( .a(N7503), .b(N10681), .O(N10746) );
nand2 gate3185( .a(N7521), .b(N10683), .O(N10747) );
nand2 gate3186( .a(N8678), .b(N10685), .O(N10748) );
nand2 gate3187( .a(N8690), .b(N10687), .O(N10749) );
nand2 gate3188( .a(N9685), .b(N10689), .O(N10750) );
nand2 gate3189( .a(N8757), .b(N10694), .O(N10753) );
nand2 gate3190( .a(N8769), .b(N10696), .O(N10754) );
or2 gate3191( .a(N10705), .b(N10549), .O(N10759) );
or2 gate3192( .a(N10707), .b(N10553), .O(N10760) );
or2 gate3193( .a(N10708), .b(N10554), .O(N10761) );
inv1 gate( .a(N10709),.O(N10709_NOT) );
inv1 gate( .a(N10555),.O(N10555_NOT));
and2 gate( .a(N10709_NOT), .b(p637), .O(EX1591) );
and2 gate( .a(N10555_NOT), .b(EX1591), .O(EX1592) );
and2 gate( .a(N10709), .b(p638), .O(EX1593) );
and2 gate( .a(N10555_NOT), .b(EX1593), .O(EX1594) );
and2 gate( .a(N10709_NOT), .b(p639), .O(EX1595) );
and2 gate( .a(N10555), .b(EX1595), .O(EX1596) );
and2 gate( .a(N10709), .b(p640), .O(EX1597) );
and2 gate( .a(N10555), .b(EX1597), .O(EX1598) );
or2  gate( .a(EX1592), .b(EX1594), .O(EX1599) );
or2  gate( .a(EX1596), .b(EX1599), .O(EX1600) );
or2  gate( .a(EX1598), .b(EX1600), .O(N10762) );
or2 gate3195( .a(N10710), .b(N10556), .O(N10763) );
nand2 gate3196( .a(N8580), .b(N10719), .O(N10764) );
and2 gate3197( .a(N10652), .b(N9890), .O(N10765) );
and2 gate3198( .a(N10652), .b(N9891), .O(N10766) );
inv1 gate( .a(N10652),.O(N10652_NOT) );
inv1 gate( .a(N9892),.O(N9892_NOT));
and2 gate( .a(N10652_NOT), .b(p641), .O(EX1601) );
and2 gate( .a(N9892_NOT), .b(EX1601), .O(EX1602) );
and2 gate( .a(N10652), .b(p642), .O(EX1603) );
and2 gate( .a(N9892_NOT), .b(EX1603), .O(EX1604) );
and2 gate( .a(N10652_NOT), .b(p643), .O(EX1605) );
and2 gate( .a(N9892), .b(EX1605), .O(EX1606) );
and2 gate( .a(N10652), .b(p644), .O(EX1607) );
and2 gate( .a(N9892), .b(EX1607), .O(EX1608) );
or2  gate( .a(EX1602), .b(EX1604), .O(EX1609) );
or2  gate( .a(EX1606), .b(EX1609), .O(EX1610) );
or2  gate( .a(EX1608), .b(EX1610), .O(N10767) );
and2 gate3200( .a(N10652), .b(N8252), .O(N10768) );
inv1 gate3201( .a(N10659), .O(N10769) );
inv1 gate( .a(N10659),.O(N10659_NOT) );
inv1 gate( .a(N9245),.O(N9245_NOT));
and2 gate( .a(N10659_NOT), .b(p645), .O(EX1611) );
and2 gate( .a(N9245_NOT), .b(EX1611), .O(EX1612) );
and2 gate( .a(N10659), .b(p646), .O(EX1613) );
and2 gate( .a(N9245_NOT), .b(EX1613), .O(EX1614) );
and2 gate( .a(N10659_NOT), .b(p647), .O(EX1615) );
and2 gate( .a(N9245), .b(EX1615), .O(EX1616) );
and2 gate( .a(N10659), .b(p648), .O(EX1617) );
and2 gate( .a(N9245), .b(EX1617), .O(EX1618) );
or2  gate( .a(EX1612), .b(EX1614), .O(EX1619) );
or2  gate( .a(EX1616), .b(EX1619), .O(EX1620) );
or2  gate( .a(EX1618), .b(EX1620), .O(N10770) );
inv1 gate3203( .a(N10662), .O(N10771) );
nand2 gate3204( .a(N10662), .b(N9246), .O(N10772) );
inv1 gate3205( .a(N10665), .O(N10773) );
nand2 gate3206( .a(N10665), .b(N9247), .O(N10774) );
inv1 gate3207( .a(N10668), .O(N10775) );
nand2 gate3208( .a(N10668), .b(N9248), .O(N10776) );
inv1 gate( .a(N10730),.O(N10730_NOT) );
inv1 gate( .a(N10587),.O(N10587_NOT));
and2 gate( .a(N10730_NOT), .b(p649), .O(EX1621) );
and2 gate( .a(N10587_NOT), .b(EX1621), .O(EX1622) );
and2 gate( .a(N10730), .b(p650), .O(EX1623) );
and2 gate( .a(N10587_NOT), .b(EX1623), .O(EX1624) );
and2 gate( .a(N10730_NOT), .b(p651), .O(EX1625) );
and2 gate( .a(N10587), .b(EX1625), .O(EX1626) );
and2 gate( .a(N10730), .b(p652), .O(EX1627) );
and2 gate( .a(N10587), .b(EX1627), .O(EX1628) );
or2  gate( .a(EX1622), .b(EX1624), .O(EX1629) );
or2  gate( .a(EX1626), .b(EX1629), .O(EX1630) );
or2  gate( .a(EX1628), .b(EX1630), .O(N10778) );
or2 gate3210( .a(N10731), .b(N10588), .O(N10781) );
inv1 gate3211( .a(N10652), .O(N10784) );
nand2 gate3212( .a(N10737), .b(N10672), .O(N10789) );
nand2 gate3213( .a(N10738), .b(N10674), .O(N10792) );
inv1 gate3214( .a(N10675), .O(N10796) );
nand2 gate3215( .a(N10675), .b(N8633), .O(N10797) );
inv1 gate3216( .a(N10678), .O(N10798) );
nand2 gate3217( .a(N10678), .b(N8638), .O(N10799) );
nand2 gate3218( .a(N10746), .b(N10682), .O(N10800) );
nand2 gate3219( .a(N10747), .b(N10684), .O(N10803) );
nand2 gate3220( .a(N10748), .b(N10686), .O(N10806) );
nand2 gate3221( .a(N10749), .b(N10688), .O(N10809) );
nand2 gate3222( .a(N10750), .b(N10690), .O(N10812) );
inv1 gate3223( .a(N10691), .O(N10815) );
nand2 gate3224( .a(N10691), .b(N9866), .O(N10816) );
inv1 gate( .a(N10753),.O(N10753_NOT) );
inv1 gate( .a(N10695),.O(N10695_NOT));
and2 gate( .a(N10753_NOT), .b(p653), .O(EX1631) );
and2 gate( .a(N10695_NOT), .b(EX1631), .O(EX1632) );
and2 gate( .a(N10753), .b(p654), .O(EX1633) );
and2 gate( .a(N10695_NOT), .b(EX1633), .O(EX1634) );
and2 gate( .a(N10753_NOT), .b(p655), .O(EX1635) );
and2 gate( .a(N10695), .b(EX1635), .O(EX1636) );
and2 gate( .a(N10753), .b(p656), .O(EX1637) );
and2 gate( .a(N10695), .b(EX1637), .O(EX1638) );
or2  gate( .a(EX1632), .b(EX1634), .O(EX1639) );
or2  gate( .a(EX1636), .b(EX1639), .O(EX1640) );
or2  gate( .a(EX1638), .b(EX1640), .O(N10817) );
nand2 gate3226( .a(N10754), .b(N10697), .O(N10820) );
inv1 gate3227( .a(N10698), .O(N10823) );
nand2 gate3228( .a(N10698), .b(N9505), .O(N10824) );
inv1 gate3229( .a(N10701), .O(N10825) );
nand2 gate3230( .a(N10701), .b(N9514), .O(N10826) );
nand2 gate3231( .a(N10764), .b(N10720), .O(N10827) );
nand2 gate3232( .a(N8583), .b(N10769), .O(N10832) );
nand2 gate3233( .a(N8586), .b(N10771), .O(N10833) );
nand2 gate3234( .a(N8589), .b(N10773), .O(N10834) );
nand2 gate3235( .a(N8592), .b(N10775), .O(N10835) );
inv1 gate3236( .a(N10739), .O(N10836) );
buf1 gate3237( .a(N10778), .O(N10837) );
buf1 gate3238( .a(N10778), .O(N10838) );
buf1 gate3239( .a(N10781), .O(N10839) );
buf1 gate3240( .a(N10781), .O(N10840) );
nand2 gate3241( .a(N7482), .b(N10796), .O(N10845) );
nand2 gate3242( .a(N7494), .b(N10798), .O(N10846) );
nand2 gate3243( .a(N9473), .b(N10815), .O(N10857) );
nand2 gate3244( .a(N8781), .b(N10823), .O(N10862) );
nand2 gate3245( .a(N8799), .b(N10825), .O(N10863) );
and2 gate3246( .a(N10023), .b(N10784), .O(N10864) );
and2 gate3247( .a(N10024), .b(N10784), .O(N10865) );
and2 gate3248( .a(N9739), .b(N10784), .O(N10866) );
inv1 gate( .a(N7136),.O(N7136_NOT) );
inv1 gate( .a(N10784),.O(N10784_NOT));
and2 gate( .a(N7136_NOT), .b(p657), .O(EX1641) );
and2 gate( .a(N10784_NOT), .b(EX1641), .O(EX1642) );
and2 gate( .a(N7136), .b(p658), .O(EX1643) );
and2 gate( .a(N10784_NOT), .b(EX1643), .O(EX1644) );
and2 gate( .a(N7136_NOT), .b(p659), .O(EX1645) );
and2 gate( .a(N10784), .b(EX1645), .O(EX1646) );
and2 gate( .a(N7136), .b(p660), .O(EX1647) );
and2 gate( .a(N10784), .b(EX1647), .O(EX1648) );
or2  gate( .a(EX1642), .b(EX1644), .O(EX1649) );
or2  gate( .a(EX1646), .b(EX1649), .O(EX1650) );
or2  gate( .a(EX1648), .b(EX1650), .O(N10867) );
nand2 gate3250( .a(N10832), .b(N10770), .O(N10868) );
nand2 gate3251( .a(N10833), .b(N10772), .O(N10869) );
nand2 gate3252( .a(N10834), .b(N10774), .O(N10870) );
nand2 gate3253( .a(N10835), .b(N10776), .O(N10871) );
inv1 gate3254( .a(N10789), .O(N10872) );
nand2 gate3255( .a(N10789), .b(N8616), .O(N10873) );
inv1 gate3256( .a(N10792), .O(N10874) );
nand2 gate3257( .a(N10792), .b(N8625), .O(N10875) );
nand2 gate3258( .a(N10845), .b(N10797), .O(N10876) );
inv1 gate( .a(N10846),.O(N10846_NOT) );
inv1 gate( .a(N10799),.O(N10799_NOT));
and2 gate( .a(N10846_NOT), .b(p661), .O(EX1651) );
and2 gate( .a(N10799_NOT), .b(EX1651), .O(EX1652) );
and2 gate( .a(N10846), .b(p662), .O(EX1653) );
and2 gate( .a(N10799_NOT), .b(EX1653), .O(EX1654) );
and2 gate( .a(N10846_NOT), .b(p663), .O(EX1655) );
and2 gate( .a(N10799), .b(EX1655), .O(EX1656) );
and2 gate( .a(N10846), .b(p664), .O(EX1657) );
and2 gate( .a(N10799), .b(EX1657), .O(EX1658) );
or2  gate( .a(EX1652), .b(EX1654), .O(EX1659) );
or2  gate( .a(EX1656), .b(EX1659), .O(EX1660) );
or2  gate( .a(EX1658), .b(EX1660), .O(N10879) );
inv1 gate3260( .a(N10800), .O(N10882) );
nand2 gate3261( .a(N10800), .b(N8645), .O(N10883) );
inv1 gate3262( .a(N10803), .O(N10884) );
inv1 gate( .a(N10803),.O(N10803_NOT) );
inv1 gate( .a(N8654),.O(N8654_NOT));
and2 gate( .a(N10803_NOT), .b(p665), .O(EX1661) );
and2 gate( .a(N8654_NOT), .b(EX1661), .O(EX1662) );
and2 gate( .a(N10803), .b(p666), .O(EX1663) );
and2 gate( .a(N8654_NOT), .b(EX1663), .O(EX1664) );
and2 gate( .a(N10803_NOT), .b(p667), .O(EX1665) );
and2 gate( .a(N8654), .b(EX1665), .O(EX1666) );
and2 gate( .a(N10803), .b(p668), .O(EX1667) );
and2 gate( .a(N8654), .b(EX1667), .O(EX1668) );
or2  gate( .a(EX1662), .b(EX1664), .O(EX1669) );
or2  gate( .a(EX1666), .b(EX1669), .O(EX1670) );
or2  gate( .a(EX1668), .b(EX1670), .O(N10885) );
inv1 gate3264( .a(N10806), .O(N10886) );
nand2 gate3265( .a(N10806), .b(N9455), .O(N10887) );
inv1 gate3266( .a(N10809), .O(N10888) );
nand2 gate3267( .a(N10809), .b(N9460), .O(N10889) );
inv1 gate3268( .a(N10812), .O(N10890) );
nand2 gate3269( .a(N10812), .b(N9862), .O(N10891) );
nand2 gate3270( .a(N10857), .b(N10816), .O(N10892) );
inv1 gate3271( .a(N10817), .O(N10895) );
nand2 gate3272( .a(N10817), .b(N9494), .O(N10896) );
inv1 gate3273( .a(N10820), .O(N10897) );
inv1 gate( .a(N10820),.O(N10820_NOT) );
inv1 gate( .a(N9499),.O(N9499_NOT));
and2 gate( .a(N10820_NOT), .b(p669), .O(EX1671) );
and2 gate( .a(N9499_NOT), .b(EX1671), .O(EX1672) );
and2 gate( .a(N10820), .b(p670), .O(EX1673) );
and2 gate( .a(N9499_NOT), .b(EX1673), .O(EX1674) );
and2 gate( .a(N10820_NOT), .b(p671), .O(EX1675) );
and2 gate( .a(N9499), .b(EX1675), .O(EX1676) );
and2 gate( .a(N10820), .b(p672), .O(EX1677) );
and2 gate( .a(N9499), .b(EX1677), .O(EX1678) );
or2  gate( .a(EX1672), .b(EX1674), .O(EX1679) );
or2  gate( .a(EX1676), .b(EX1679), .O(EX1680) );
or2  gate( .a(EX1678), .b(EX1680), .O(N10898) );
nand2 gate3275( .a(N10862), .b(N10824), .O(N10899) );
nand2 gate3276( .a(N10863), .b(N10826), .O(N10902) );
or2 gate3277( .a(N10864), .b(N10765), .O(N10905) );
or2 gate3278( .a(N10865), .b(N10766), .O(N10906) );
or2 gate3279( .a(N10866), .b(N10767), .O(N10907) );
or2 gate3280( .a(N10867), .b(N10768), .O(N10908) );
nand2 gate3281( .a(N7450), .b(N10872), .O(N10909) );
nand2 gate3282( .a(N7468), .b(N10874), .O(N10910) );
nand2 gate3283( .a(N7506), .b(N10882), .O(N10915) );
nand2 gate3284( .a(N7524), .b(N10884), .O(N10916) );
inv1 gate( .a(N8681),.O(N8681_NOT) );
inv1 gate( .a(N10886),.O(N10886_NOT));
and2 gate( .a(N8681_NOT), .b(p673), .O(EX1681) );
and2 gate( .a(N10886_NOT), .b(EX1681), .O(EX1682) );
and2 gate( .a(N8681), .b(p674), .O(EX1683) );
and2 gate( .a(N10886_NOT), .b(EX1683), .O(EX1684) );
and2 gate( .a(N8681_NOT), .b(p675), .O(EX1685) );
and2 gate( .a(N10886), .b(EX1685), .O(EX1686) );
and2 gate( .a(N8681), .b(p676), .O(EX1687) );
and2 gate( .a(N10886), .b(EX1687), .O(EX1688) );
or2  gate( .a(EX1682), .b(EX1684), .O(EX1689) );
or2  gate( .a(EX1686), .b(EX1689), .O(EX1690) );
or2  gate( .a(EX1688), .b(EX1690), .O(N10917) );
nand2 gate3286( .a(N8693), .b(N10888), .O(N10918) );
nand2 gate3287( .a(N9462), .b(N10890), .O(N10919) );
nand2 gate3288( .a(N8760), .b(N10895), .O(N10922) );
nand2 gate3289( .a(N8772), .b(N10897), .O(N10923) );
nand2 gate3290( .a(N10909), .b(N10873), .O(N10928) );
nand2 gate3291( .a(N10910), .b(N10875), .O(N10931) );
inv1 gate3292( .a(N10876), .O(N10934) );
inv1 gate( .a(N10876),.O(N10876_NOT) );
inv1 gate( .a(N8634),.O(N8634_NOT));
and2 gate( .a(N10876_NOT), .b(p677), .O(EX1691) );
and2 gate( .a(N8634_NOT), .b(EX1691), .O(EX1692) );
and2 gate( .a(N10876), .b(p678), .O(EX1693) );
and2 gate( .a(N8634_NOT), .b(EX1693), .O(EX1694) );
and2 gate( .a(N10876_NOT), .b(p679), .O(EX1695) );
and2 gate( .a(N8634), .b(EX1695), .O(EX1696) );
and2 gate( .a(N10876), .b(p680), .O(EX1697) );
and2 gate( .a(N8634), .b(EX1697), .O(EX1698) );
or2  gate( .a(EX1692), .b(EX1694), .O(EX1699) );
or2  gate( .a(EX1696), .b(EX1699), .O(EX1700) );
or2  gate( .a(EX1698), .b(EX1700), .O(N10935) );
inv1 gate3294( .a(N10879), .O(N10936) );
nand2 gate3295( .a(N10879), .b(N8639), .O(N10937) );
nand2 gate3296( .a(N10915), .b(N10883), .O(N10938) );
nand2 gate3297( .a(N10916), .b(N10885), .O(N10941) );
inv1 gate( .a(N10917),.O(N10917_NOT) );
inv1 gate( .a(N10887),.O(N10887_NOT));
and2 gate( .a(N10917_NOT), .b(p681), .O(EX1701) );
and2 gate( .a(N10887_NOT), .b(EX1701), .O(EX1702) );
and2 gate( .a(N10917), .b(p682), .O(EX1703) );
and2 gate( .a(N10887_NOT), .b(EX1703), .O(EX1704) );
and2 gate( .a(N10917_NOT), .b(p683), .O(EX1705) );
and2 gate( .a(N10887), .b(EX1705), .O(EX1706) );
and2 gate( .a(N10917), .b(p684), .O(EX1707) );
and2 gate( .a(N10887), .b(EX1707), .O(EX1708) );
or2  gate( .a(EX1702), .b(EX1704), .O(EX1709) );
or2  gate( .a(EX1706), .b(EX1709), .O(EX1710) );
or2  gate( .a(EX1708), .b(EX1710), .O(N10944) );
nand2 gate3299( .a(N10918), .b(N10889), .O(N10947) );
nand2 gate3300( .a(N10919), .b(N10891), .O(N10950) );
inv1 gate3301( .a(N10892), .O(N10953) );
nand2 gate3302( .a(N10892), .b(N9476), .O(N10954) );
nand2 gate3303( .a(N10922), .b(N10896), .O(N10955) );
nand2 gate3304( .a(N10923), .b(N10898), .O(N10958) );
inv1 gate3305( .a(N10899), .O(N10961) );
nand2 gate3306( .a(N10899), .b(N9506), .O(N10962) );
inv1 gate3307( .a(N10902), .O(N10963) );
nand2 gate3308( .a(N10902), .b(N9515), .O(N10964) );
nand2 gate3309( .a(N7485), .b(N10934), .O(N10969) );
nand2 gate3310( .a(N7497), .b(N10936), .O(N10970) );
nand2 gate3311( .a(N8718), .b(N10953), .O(N10981) );
nand2 gate3312( .a(N8784), .b(N10961), .O(N10986) );
nand2 gate3313( .a(N8802), .b(N10963), .O(N10987) );
inv1 gate3314( .a(N10928), .O(N10988) );
nand2 gate3315( .a(N10928), .b(N8617), .O(N10989) );
inv1 gate3316( .a(N10931), .O(N10990) );
nand2 gate3317( .a(N10931), .b(N8626), .O(N10991) );
nand2 gate3318( .a(N10969), .b(N10935), .O(N10992) );
nand2 gate3319( .a(N10970), .b(N10937), .O(N10995) );
inv1 gate3320( .a(N10938), .O(N10998) );
nand2 gate3321( .a(N10938), .b(N8646), .O(N10999) );
inv1 gate3322( .a(N10941), .O(N11000) );
nand2 gate3323( .a(N10941), .b(N8655), .O(N11001) );
inv1 gate3324( .a(N10944), .O(N11002) );
nand2 gate3325( .a(N10944), .b(N9456), .O(N11003) );
inv1 gate3326( .a(N10947), .O(N11004) );
nand2 gate3327( .a(N10947), .b(N9461), .O(N11005) );
inv1 gate3328( .a(N10950), .O(N11006) );
nand2 gate3329( .a(N10950), .b(N9465), .O(N11007) );
nand2 gate3330( .a(N10981), .b(N10954), .O(N11008) );
inv1 gate3331( .a(N10955), .O(N11011) );
nand2 gate3332( .a(N10955), .b(N9495), .O(N11012) );
inv1 gate3333( .a(N10958), .O(N11013) );
nand2 gate3334( .a(N10958), .b(N9500), .O(N11014) );
nand2 gate3335( .a(N10986), .b(N10962), .O(N11015) );
nand2 gate3336( .a(N10987), .b(N10964), .O(N11018) );
nand2 gate3337( .a(N7453), .b(N10988), .O(N11023) );
nand2 gate3338( .a(N7471), .b(N10990), .O(N11024) );
nand2 gate3339( .a(N7509), .b(N10998), .O(N11027) );
nand2 gate3340( .a(N7527), .b(N11000), .O(N11028) );
nand2 gate3341( .a(N8684), .b(N11002), .O(N11029) );
nand2 gate3342( .a(N8696), .b(N11004), .O(N11030) );
nand2 gate3343( .a(N8702), .b(N11006), .O(N11031) );
nand2 gate3344( .a(N8763), .b(N11011), .O(N11034) );
nand2 gate3345( .a(N8775), .b(N11013), .O(N11035) );
inv1 gate3346( .a(N10992), .O(N11040) );
nand2 gate3347( .a(N10992), .b(N8294), .O(N11041) );
inv1 gate3348( .a(N10995), .O(N11042) );
nand2 gate3349( .a(N10995), .b(N8295), .O(N11043) );
nand2 gate3350( .a(N11023), .b(N10989), .O(N11044) );
nand2 gate3351( .a(N11024), .b(N10991), .O(N11047) );
nand2 gate3352( .a(N11027), .b(N10999), .O(N11050) );
nand2 gate3353( .a(N11028), .b(N11001), .O(N11053) );
inv1 gate( .a(N11029),.O(N11029_NOT) );
inv1 gate( .a(N11003),.O(N11003_NOT));
and2 gate( .a(N11029_NOT), .b(p685), .O(EX1711) );
and2 gate( .a(N11003_NOT), .b(EX1711), .O(EX1712) );
and2 gate( .a(N11029), .b(p686), .O(EX1713) );
and2 gate( .a(N11003_NOT), .b(EX1713), .O(EX1714) );
and2 gate( .a(N11029_NOT), .b(p687), .O(EX1715) );
and2 gate( .a(N11003), .b(EX1715), .O(EX1716) );
and2 gate( .a(N11029), .b(p688), .O(EX1717) );
and2 gate( .a(N11003), .b(EX1717), .O(EX1718) );
or2  gate( .a(EX1712), .b(EX1714), .O(EX1719) );
or2  gate( .a(EX1716), .b(EX1719), .O(EX1720) );
or2  gate( .a(EX1718), .b(EX1720), .O(N11056) );
nand2 gate3355( .a(N11030), .b(N11005), .O(N11059) );
nand2 gate3356( .a(N11031), .b(N11007), .O(N11062) );
inv1 gate3357( .a(N11008), .O(N11065) );
nand2 gate3358( .a(N11008), .b(N9477), .O(N11066) );
nand2 gate3359( .a(N11034), .b(N11012), .O(N11067) );
nand2 gate3360( .a(N11035), .b(N11014), .O(N11070) );
inv1 gate3361( .a(N11015), .O(N11073) );
nand2 gate3362( .a(N11015), .b(N9507), .O(N11074) );
inv1 gate3363( .a(N11018), .O(N11075) );
nand2 gate3364( .a(N11018), .b(N9516), .O(N11076) );
nand2 gate3365( .a(N7488), .b(N11040), .O(N11077) );
inv1 gate( .a(N7500),.O(N7500_NOT) );
inv1 gate( .a(N11042),.O(N11042_NOT));
and2 gate( .a(N7500_NOT), .b(p689), .O(EX1721) );
and2 gate( .a(N11042_NOT), .b(EX1721), .O(EX1722) );
and2 gate( .a(N7500), .b(p690), .O(EX1723) );
and2 gate( .a(N11042_NOT), .b(EX1723), .O(EX1724) );
and2 gate( .a(N7500_NOT), .b(p691), .O(EX1725) );
and2 gate( .a(N11042), .b(EX1725), .O(EX1726) );
and2 gate( .a(N7500), .b(p692), .O(EX1727) );
and2 gate( .a(N11042), .b(EX1727), .O(EX1728) );
or2  gate( .a(EX1722), .b(EX1724), .O(EX1729) );
or2  gate( .a(EX1726), .b(EX1729), .O(EX1730) );
or2  gate( .a(EX1728), .b(EX1730), .O(N11078) );
nand2 gate3367( .a(N8721), .b(N11065), .O(N11095) );
nand2 gate3368( .a(N8787), .b(N11073), .O(N11098) );
inv1 gate( .a(N8805),.O(N8805_NOT) );
inv1 gate( .a(N11075),.O(N11075_NOT));
and2 gate( .a(N8805_NOT), .b(p693), .O(EX1731) );
and2 gate( .a(N11075_NOT), .b(EX1731), .O(EX1732) );
and2 gate( .a(N8805), .b(p694), .O(EX1733) );
and2 gate( .a(N11075_NOT), .b(EX1733), .O(EX1734) );
and2 gate( .a(N8805_NOT), .b(p695), .O(EX1735) );
and2 gate( .a(N11075), .b(EX1735), .O(EX1736) );
and2 gate( .a(N8805), .b(p696), .O(EX1737) );
and2 gate( .a(N11075), .b(EX1737), .O(EX1738) );
or2  gate( .a(EX1732), .b(EX1734), .O(EX1739) );
or2  gate( .a(EX1736), .b(EX1739), .O(EX1740) );
or2  gate( .a(EX1738), .b(EX1740), .O(N11099) );
nand2 gate3370( .a(N11077), .b(N11041), .O(N11100) );
nand2 gate3371( .a(N11078), .b(N11043), .O(N11103) );
inv1 gate3372( .a(N11056), .O(N11106) );
inv1 gate( .a(N11056),.O(N11056_NOT) );
inv1 gate( .a(N9319),.O(N9319_NOT));
and2 gate( .a(N11056_NOT), .b(p697), .O(EX1741) );
and2 gate( .a(N9319_NOT), .b(EX1741), .O(EX1742) );
and2 gate( .a(N11056), .b(p698), .O(EX1743) );
and2 gate( .a(N9319_NOT), .b(EX1743), .O(EX1744) );
and2 gate( .a(N11056_NOT), .b(p699), .O(EX1745) );
and2 gate( .a(N9319), .b(EX1745), .O(EX1746) );
and2 gate( .a(N11056), .b(p700), .O(EX1747) );
and2 gate( .a(N9319), .b(EX1747), .O(EX1748) );
or2  gate( .a(EX1742), .b(EX1744), .O(EX1749) );
or2  gate( .a(EX1746), .b(EX1749), .O(EX1750) );
or2  gate( .a(EX1748), .b(EX1750), .O(N11107) );
inv1 gate3374( .a(N11059), .O(N11108) );
nand2 gate3375( .a(N11059), .b(N9320), .O(N11109) );
inv1 gate3376( .a(N11067), .O(N11110) );
nand2 gate3377( .a(N11067), .b(N9381), .O(N11111) );
inv1 gate3378( .a(N11070), .O(N11112) );
nand2 gate3379( .a(N11070), .b(N9382), .O(N11113) );
inv1 gate3380( .a(N11044), .O(N11114) );
nand2 gate3381( .a(N11044), .b(N8618), .O(N11115) );
inv1 gate3382( .a(N11047), .O(N11116) );
nand2 gate3383( .a(N11047), .b(N8619), .O(N11117) );
inv1 gate3384( .a(N11050), .O(N11118) );
nand2 gate3385( .a(N11050), .b(N8647), .O(N11119) );
inv1 gate3386( .a(N11053), .O(N11120) );
nand2 gate3387( .a(N11053), .b(N8648), .O(N11121) );
inv1 gate3388( .a(N11062), .O(N11122) );
nand2 gate3389( .a(N11062), .b(N9466), .O(N11123) );
nand2 gate3390( .a(N11095), .b(N11066), .O(N11124) );
nand2 gate3391( .a(N11098), .b(N11074), .O(N11127) );
nand2 gate3392( .a(N11099), .b(N11076), .O(N11130) );
nand2 gate3393( .a(N8687), .b(N11106), .O(N11137) );
nand2 gate3394( .a(N8699), .b(N11108), .O(N11138) );
nand2 gate3395( .a(N8766), .b(N11110), .O(N11139) );
inv1 gate( .a(N8778),.O(N8778_NOT) );
inv1 gate( .a(N11112),.O(N11112_NOT));
and2 gate( .a(N8778_NOT), .b(p701), .O(EX1751) );
and2 gate( .a(N11112_NOT), .b(EX1751), .O(EX1752) );
and2 gate( .a(N8778), .b(p702), .O(EX1753) );
and2 gate( .a(N11112_NOT), .b(EX1753), .O(EX1754) );
and2 gate( .a(N8778_NOT), .b(p703), .O(EX1755) );
and2 gate( .a(N11112), .b(EX1755), .O(EX1756) );
and2 gate( .a(N8778), .b(p704), .O(EX1757) );
and2 gate( .a(N11112), .b(EX1757), .O(EX1758) );
or2  gate( .a(EX1752), .b(EX1754), .O(EX1759) );
or2  gate( .a(EX1756), .b(EX1759), .O(EX1760) );
or2  gate( .a(EX1758), .b(EX1760), .O(N11140) );
nand2 gate3397( .a(N7456), .b(N11114), .O(N11141) );
nand2 gate3398( .a(N7474), .b(N11116), .O(N11142) );
inv1 gate( .a(N7512),.O(N7512_NOT) );
inv1 gate( .a(N11118),.O(N11118_NOT));
and2 gate( .a(N7512_NOT), .b(p705), .O(EX1761) );
and2 gate( .a(N11118_NOT), .b(EX1761), .O(EX1762) );
and2 gate( .a(N7512), .b(p706), .O(EX1763) );
and2 gate( .a(N11118_NOT), .b(EX1763), .O(EX1764) );
and2 gate( .a(N7512_NOT), .b(p707), .O(EX1765) );
and2 gate( .a(N11118), .b(EX1765), .O(EX1766) );
and2 gate( .a(N7512), .b(p708), .O(EX1767) );
and2 gate( .a(N11118), .b(EX1767), .O(EX1768) );
or2  gate( .a(EX1762), .b(EX1764), .O(EX1769) );
or2  gate( .a(EX1766), .b(EX1769), .O(EX1770) );
or2  gate( .a(EX1768), .b(EX1770), .O(N11143) );
nand2 gate3400( .a(N7530), .b(N11120), .O(N11144) );
inv1 gate( .a(N8705),.O(N8705_NOT) );
inv1 gate( .a(N11122),.O(N11122_NOT));
and2 gate( .a(N8705_NOT), .b(p709), .O(EX1771) );
and2 gate( .a(N11122_NOT), .b(EX1771), .O(EX1772) );
and2 gate( .a(N8705), .b(p710), .O(EX1773) );
and2 gate( .a(N11122_NOT), .b(EX1773), .O(EX1774) );
and2 gate( .a(N8705_NOT), .b(p711), .O(EX1775) );
and2 gate( .a(N11122), .b(EX1775), .O(EX1776) );
and2 gate( .a(N8705), .b(p712), .O(EX1777) );
and2 gate( .a(N11122), .b(EX1777), .O(EX1778) );
or2  gate( .a(EX1772), .b(EX1774), .O(EX1779) );
or2  gate( .a(EX1776), .b(EX1779), .O(EX1780) );
or2  gate( .a(EX1778), .b(EX1780), .O(N11145) );
and3 gate3402( .a(N11103), .b(N8871), .c(N10283), .O(N11152) );
and3 gate3403( .a(N11100), .b(N7655), .c(N10283), .O(N11153) );
and3 gate3404( .a(N11103), .b(N9551), .c(N10119), .O(N11154) );
and3 gate3405( .a(N11100), .b(N9917), .c(N10119), .O(N11155) );
nand2 gate3406( .a(N11137), .b(N11107), .O(N11156) );
nand2 gate3407( .a(N11138), .b(N11109), .O(N11159) );
nand2 gate3408( .a(N11139), .b(N11111), .O(N11162) );
nand2 gate3409( .a(N11140), .b(N11113), .O(N11165) );
nand2 gate3410( .a(N11141), .b(N11115), .O(N11168) );
nand2 gate3411( .a(N11142), .b(N11117), .O(N11171) );
nand2 gate3412( .a(N11143), .b(N11119), .O(N11174) );
nand2 gate3413( .a(N11144), .b(N11121), .O(N11177) );
nand2 gate3414( .a(N11145), .b(N11123), .O(N11180) );
inv1 gate3415( .a(N11124), .O(N11183) );
nand2 gate3416( .a(N11124), .b(N9468), .O(N11184) );
inv1 gate3417( .a(N11127), .O(N11185) );
nand2 gate3418( .a(N11127), .b(N9508), .O(N11186) );
inv1 gate3419( .a(N11130), .O(N11187) );
inv1 gate( .a(N11130),.O(N11130_NOT) );
inv1 gate( .a(N9509),.O(N9509_NOT));
and2 gate( .a(N11130_NOT), .b(p713), .O(EX1781) );
and2 gate( .a(N9509_NOT), .b(EX1781), .O(EX1782) );
and2 gate( .a(N11130), .b(p714), .O(EX1783) );
and2 gate( .a(N9509_NOT), .b(EX1783), .O(EX1784) );
and2 gate( .a(N11130_NOT), .b(p715), .O(EX1785) );
and2 gate( .a(N9509), .b(EX1785), .O(EX1786) );
and2 gate( .a(N11130), .b(p716), .O(EX1787) );
and2 gate( .a(N9509), .b(EX1787), .O(EX1788) );
or2  gate( .a(EX1782), .b(EX1784), .O(EX1789) );
or2  gate( .a(EX1786), .b(EX1789), .O(EX1790) );
or2  gate( .a(EX1788), .b(EX1790), .O(N11188) );
or4 gate3421( .a(N11152), .b(N11153), .c(N11154), .d(N11155), .O(N11205) );
nand2 gate3422( .a(N8724), .b(N11183), .O(N11210) );
inv1 gate( .a(N8790),.O(N8790_NOT) );
inv1 gate( .a(N11185),.O(N11185_NOT));
and2 gate( .a(N8790_NOT), .b(p717), .O(EX1791) );
and2 gate( .a(N11185_NOT), .b(EX1791), .O(EX1792) );
and2 gate( .a(N8790), .b(p718), .O(EX1793) );
and2 gate( .a(N11185_NOT), .b(EX1793), .O(EX1794) );
and2 gate( .a(N8790_NOT), .b(p719), .O(EX1795) );
and2 gate( .a(N11185), .b(EX1795), .O(EX1796) );
and2 gate( .a(N8790), .b(p720), .O(EX1797) );
and2 gate( .a(N11185), .b(EX1797), .O(EX1798) );
or2  gate( .a(EX1792), .b(EX1794), .O(EX1799) );
or2  gate( .a(EX1796), .b(EX1799), .O(EX1800) );
or2  gate( .a(EX1798), .b(EX1800), .O(N11211) );
nand2 gate3424( .a(N8808), .b(N11187), .O(N11212) );
inv1 gate3425( .a(N11168), .O(N11213) );
nand2 gate3426( .a(N11168), .b(N8260), .O(N11214) );
inv1 gate3427( .a(N11171), .O(N11215) );
nand2 gate3428( .a(N11171), .b(N8261), .O(N11216) );
inv1 gate3429( .a(N11174), .O(N11217) );
nand2 gate3430( .a(N11174), .b(N8296), .O(N11218) );
inv1 gate3431( .a(N11177), .O(N11219) );
nand2 gate3432( .a(N11177), .b(N8297), .O(N11220) );
and3 gate3433( .a(N11159), .b(N9575), .c(N1218), .O(N11222) );
and3 gate3434( .a(N11156), .b(N8927), .c(N1218), .O(N11223) );
and3 gate3435( .a(N11159), .b(N9935), .c(N750), .O(N11224) );
and3 gate3436( .a(N11156), .b(N10132), .c(N750), .O(N11225) );
and3 gate3437( .a(N11165), .b(N9608), .c(N10497), .O(N11226) );
and3 gate3438( .a(N11162), .b(N9001), .c(N10497), .O(N11227) );
and3 gate3439( .a(N11165), .b(N9949), .c(N10301), .O(N11228) );
and3 gate3440( .a(N11162), .b(N10160), .c(N10301), .O(N11229) );
inv1 gate3441( .a(N11180), .O(N11231) );
nand2 gate3442( .a(N11180), .b(N9467), .O(N11232) );
nand2 gate3443( .a(N11210), .b(N11184), .O(N11233) );
nand2 gate3444( .a(N11211), .b(N11186), .O(N11236) );
nand2 gate3445( .a(N11212), .b(N11188), .O(N11239) );
nand2 gate3446( .a(N7459), .b(N11213), .O(N11242) );
inv1 gate( .a(N7462),.O(N7462_NOT) );
inv1 gate( .a(N11215),.O(N11215_NOT));
and2 gate( .a(N7462_NOT), .b(p721), .O(EX1801) );
and2 gate( .a(N11215_NOT), .b(EX1801), .O(EX1802) );
and2 gate( .a(N7462), .b(p722), .O(EX1803) );
and2 gate( .a(N11215_NOT), .b(EX1803), .O(EX1804) );
and2 gate( .a(N7462_NOT), .b(p723), .O(EX1805) );
and2 gate( .a(N11215), .b(EX1805), .O(EX1806) );
and2 gate( .a(N7462), .b(p724), .O(EX1807) );
and2 gate( .a(N11215), .b(EX1807), .O(EX1808) );
or2  gate( .a(EX1802), .b(EX1804), .O(EX1809) );
or2  gate( .a(EX1806), .b(EX1809), .O(EX1810) );
or2  gate( .a(EX1808), .b(EX1810), .O(N11243) );
nand2 gate3448( .a(N7515), .b(N11217), .O(N11244) );
nand2 gate3449( .a(N7518), .b(N11219), .O(N11245) );
inv1 gate3450( .a(N11205), .O(N11246) );
nand2 gate3451( .a(N8708), .b(N11231), .O(N11250) );
or4 gate3452( .a(N11222), .b(N11223), .c(N11224), .d(N11225), .O(N11252) );
or4 gate3453( .a(N11226), .b(N11227), .c(N11228), .d(N11229), .O(N11257) );
nand2 gate3454( .a(N11242), .b(N11214), .O(N11260) );
nand2 gate3455( .a(N11243), .b(N11216), .O(N11261) );
nand2 gate3456( .a(N11244), .b(N11218), .O(N11262) );
nand2 gate3457( .a(N11245), .b(N11220), .O(N11263) );
inv1 gate3458( .a(N11233), .O(N11264) );
nand2 gate3459( .a(N11233), .b(N9322), .O(N11265) );
inv1 gate3460( .a(N11236), .O(N11267) );
inv1 gate( .a(N11236),.O(N11236_NOT) );
inv1 gate( .a(N9383),.O(N9383_NOT));
and2 gate( .a(N11236_NOT), .b(p725), .O(EX1811) );
and2 gate( .a(N9383_NOT), .b(EX1811), .O(EX1812) );
and2 gate( .a(N11236), .b(p726), .O(EX1813) );
and2 gate( .a(N9383_NOT), .b(EX1813), .O(EX1814) );
and2 gate( .a(N11236_NOT), .b(p727), .O(EX1815) );
and2 gate( .a(N9383), .b(EX1815), .O(EX1816) );
and2 gate( .a(N11236), .b(p728), .O(EX1817) );
and2 gate( .a(N9383), .b(EX1817), .O(EX1818) );
or2  gate( .a(EX1812), .b(EX1814), .O(EX1819) );
or2  gate( .a(EX1816), .b(EX1819), .O(EX1820) );
or2  gate( .a(EX1818), .b(EX1820), .O(N11268) );
inv1 gate3462( .a(N11239), .O(N11269) );
nand2 gate3463( .a(N11239), .b(N9384), .O(N11270) );
nand2 gate3464( .a(N11250), .b(N11232), .O(N11272) );
inv1 gate3465( .a(N11261), .O(N11277) );
and2 gate3466( .a(N10273), .b(N11260), .O(N11278) );
inv1 gate3467( .a(N11263), .O(N11279) );
and2 gate3468( .a(N10119), .b(N11262), .O(N11280) );
nand2 gate3469( .a(N8714), .b(N11264), .O(N11282) );
inv1 gate3470( .a(N11252), .O(N11283) );
nand2 gate3471( .a(N8793), .b(N11267), .O(N11284) );
inv1 gate( .a(N8796),.O(N8796_NOT) );
inv1 gate( .a(N11269),.O(N11269_NOT));
and2 gate( .a(N8796_NOT), .b(p729), .O(EX1821) );
and2 gate( .a(N11269_NOT), .b(EX1821), .O(EX1822) );
and2 gate( .a(N8796), .b(p730), .O(EX1823) );
and2 gate( .a(N11269_NOT), .b(EX1823), .O(EX1824) );
and2 gate( .a(N8796_NOT), .b(p731), .O(EX1825) );
and2 gate( .a(N11269), .b(EX1825), .O(EX1826) );
and2 gate( .a(N8796), .b(p732), .O(EX1827) );
and2 gate( .a(N11269), .b(EX1827), .O(EX1828) );
or2  gate( .a(EX1822), .b(EX1824), .O(EX1829) );
or2  gate( .a(EX1826), .b(EX1829), .O(EX1830) );
or2  gate( .a(EX1828), .b(EX1830), .O(N11285) );
inv1 gate3473( .a(N11257), .O(N11286) );
and2 gate3474( .a(N11277), .b(N10479), .O(N11288) );
inv1 gate( .a(N11279),.O(N11279_NOT) );
inv1 gate( .a(N10283),.O(N10283_NOT));
and2 gate( .a(N11279_NOT), .b(p733), .O(EX1831) );
and2 gate( .a(N10283_NOT), .b(EX1831), .O(EX1832) );
and2 gate( .a(N11279), .b(p734), .O(EX1833) );
and2 gate( .a(N10283_NOT), .b(EX1833), .O(EX1834) );
and2 gate( .a(N11279_NOT), .b(p735), .O(EX1835) );
and2 gate( .a(N10283), .b(EX1835), .O(EX1836) );
and2 gate( .a(N11279), .b(p736), .O(EX1837) );
and2 gate( .a(N10283), .b(EX1837), .O(EX1838) );
or2  gate( .a(EX1832), .b(EX1834), .O(EX1839) );
or2  gate( .a(EX1836), .b(EX1839), .O(EX1840) );
or2  gate( .a(EX1838), .b(EX1840), .O(N11289) );
inv1 gate3476( .a(N11272), .O(N11290) );
inv1 gate( .a(N11272),.O(N11272_NOT) );
inv1 gate( .a(N9321),.O(N9321_NOT));
and2 gate( .a(N11272_NOT), .b(p737), .O(EX1841) );
and2 gate( .a(N9321_NOT), .b(EX1841), .O(EX1842) );
and2 gate( .a(N11272), .b(p738), .O(EX1843) );
and2 gate( .a(N9321_NOT), .b(EX1843), .O(EX1844) );
and2 gate( .a(N11272_NOT), .b(p739), .O(EX1845) );
and2 gate( .a(N9321), .b(EX1845), .O(EX1846) );
and2 gate( .a(N11272), .b(p740), .O(EX1847) );
and2 gate( .a(N9321), .b(EX1847), .O(EX1848) );
or2  gate( .a(EX1842), .b(EX1844), .O(EX1849) );
or2  gate( .a(EX1846), .b(EX1849), .O(EX1850) );
or2  gate( .a(EX1848), .b(EX1850), .O(N11291) );
inv1 gate( .a(N11282),.O(N11282_NOT) );
inv1 gate( .a(N11265),.O(N11265_NOT));
and2 gate( .a(N11282_NOT), .b(p741), .O(EX1851) );
and2 gate( .a(N11265_NOT), .b(EX1851), .O(EX1852) );
and2 gate( .a(N11282), .b(p742), .O(EX1853) );
and2 gate( .a(N11265_NOT), .b(EX1853), .O(EX1854) );
and2 gate( .a(N11282_NOT), .b(p743), .O(EX1855) );
and2 gate( .a(N11265), .b(EX1855), .O(EX1856) );
and2 gate( .a(N11282), .b(p744), .O(EX1857) );
and2 gate( .a(N11265), .b(EX1857), .O(EX1858) );
or2  gate( .a(EX1852), .b(EX1854), .O(EX1859) );
or2  gate( .a(EX1856), .b(EX1859), .O(EX1860) );
or2  gate( .a(EX1858), .b(EX1860), .O(N11292) );
nand2 gate3479( .a(N11284), .b(N11268), .O(N11293) );
nand2 gate3480( .a(N11285), .b(N11270), .O(N11294) );
nand2 gate3481( .a(N8711), .b(N11290), .O(N11295) );
inv1 gate3482( .a(N11292), .O(N11296) );
inv1 gate3483( .a(N11294), .O(N11297) );
and2 gate3484( .a(N10301), .b(N11293), .O(N11298) );
or2 gate3485( .a(N11288), .b(N11278), .O(N11299) );
or2 gate3486( .a(N11289), .b(N11280), .O(N11302) );
nand2 gate3487( .a(N11295), .b(N11291), .O(N11307) );
and2 gate3488( .a(N11296), .b(N1218), .O(N11308) );
and2 gate3489( .a(N11297), .b(N10497), .O(N11309) );
nand2 gate3490( .a(N11302), .b(N11246), .O(N11312) );
nand2 gate3491( .a(N11299), .b(N10836), .O(N11313) );
inv1 gate3492( .a(N11299), .O(N11314) );
inv1 gate3493( .a(N11302), .O(N11315) );
and2 gate3494( .a(N750), .b(N11307), .O(N11316) );
or2 gate3495( .a(N11309), .b(N11298), .O(N11317) );
nand2 gate3496( .a(N11205), .b(N11315), .O(N11320) );
nand2 gate3497( .a(N10739), .b(N11314), .O(N11321) );
or2 gate3498( .a(N11308), .b(N11316), .O(N11323) );
inv1 gate( .a(N11312),.O(N11312_NOT) );
inv1 gate( .a(N11320),.O(N11320_NOT));
and2 gate( .a(N11312_NOT), .b(p745), .O(EX1861) );
and2 gate( .a(N11320_NOT), .b(EX1861), .O(EX1862) );
and2 gate( .a(N11312), .b(p746), .O(EX1863) );
and2 gate( .a(N11320_NOT), .b(EX1863), .O(EX1864) );
and2 gate( .a(N11312_NOT), .b(p747), .O(EX1865) );
and2 gate( .a(N11320), .b(EX1865), .O(EX1866) );
and2 gate( .a(N11312), .b(p748), .O(EX1867) );
and2 gate( .a(N11320), .b(EX1867), .O(EX1868) );
or2  gate( .a(EX1862), .b(EX1864), .O(EX1869) );
or2  gate( .a(EX1866), .b(EX1869), .O(EX1870) );
or2  gate( .a(EX1868), .b(EX1870), .O(N11327) );
inv1 gate( .a(N11313),.O(N11313_NOT) );
inv1 gate( .a(N11321),.O(N11321_NOT));
and2 gate( .a(N11313_NOT), .b(p749), .O(EX1871) );
and2 gate( .a(N11321_NOT), .b(EX1871), .O(EX1872) );
and2 gate( .a(N11313), .b(p750), .O(EX1873) );
and2 gate( .a(N11321_NOT), .b(EX1873), .O(EX1874) );
and2 gate( .a(N11313_NOT), .b(p751), .O(EX1875) );
and2 gate( .a(N11321), .b(EX1875), .O(EX1876) );
and2 gate( .a(N11313), .b(p752), .O(EX1877) );
and2 gate( .a(N11321), .b(EX1877), .O(EX1878) );
or2  gate( .a(EX1872), .b(EX1874), .O(EX1879) );
or2  gate( .a(EX1876), .b(EX1879), .O(EX1880) );
or2  gate( .a(EX1878), .b(EX1880), .O(N11328) );
inv1 gate( .a(N11317),.O(N11317_NOT) );
inv1 gate( .a(N11286),.O(N11286_NOT));
and2 gate( .a(N11317_NOT), .b(p753), .O(EX1881) );
and2 gate( .a(N11286_NOT), .b(EX1881), .O(EX1882) );
and2 gate( .a(N11317), .b(p754), .O(EX1883) );
and2 gate( .a(N11286_NOT), .b(EX1883), .O(EX1884) );
and2 gate( .a(N11317_NOT), .b(p755), .O(EX1885) );
and2 gate( .a(N11286), .b(EX1885), .O(EX1886) );
and2 gate( .a(N11317), .b(p756), .O(EX1887) );
and2 gate( .a(N11286), .b(EX1887), .O(EX1888) );
or2  gate( .a(EX1882), .b(EX1884), .O(EX1889) );
or2  gate( .a(EX1886), .b(EX1889), .O(EX1890) );
or2  gate( .a(EX1888), .b(EX1890), .O(N11329) );
inv1 gate3502( .a(N11317), .O(N11331) );
inv1 gate3503( .a(N11327), .O(N11333) );
inv1 gate3504( .a(N11328), .O(N11334) );
nand2 gate3505( .a(N11257), .b(N11331), .O(N11335) );
nand2 gate3506( .a(N11323), .b(N11283), .O(N11336) );
inv1 gate3507( .a(N11323), .O(N11337) );
nand2 gate3508( .a(N11329), .b(N11335), .O(N11338) );
nand2 gate3509( .a(N11252), .b(N11337), .O(N11339) );
inv1 gate3510( .a(N11338), .O(N11340) );
nand2 gate3511( .a(N11336), .b(N11339), .O(N11341) );
inv1 gate3512( .a(N11341), .O(N11342) );
buf1 gate3513( .a(N241_I), .O(N241_O) );

endmodule
